// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:00 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UXrHYSFFatkkhfkDxDViu3cfxdzsTPfKStN0gI68QpV73DD/ZEK+1COuRknyY/gg
sToA22Toe88ee7FmS/m8BkTWi4Xaitw/TpcJ6bDVCtO+KPxYfkyrMAyFQTpEgy3V
5YvBR0WJvFrELPDl5tIwlJXPyqByU87rRCEVC2Q5frg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8304)
GLbpznGF00GXB+M9Gqo7LG6ZpnECgz0dF2YVGqspbS9MGgWjSkmicr2Fqn9M6a50
P4/oUDmAcaDuSXIIL7r82EMY26b9bW/EdUeIemyBu4WfiERMGuGpeBTi5zHL0DTp
5CPPTmCUDBChl9xhxwgw9sTg92DKGqw24SDRYItD3a6MP1IUYtIkSr42Twz199W7
vj8c45Ubpb7koJ8tcRyaas5uaTucRHwYBWoxItY5SkNMpILxMzFo29zvLA0y3Yvf
DR5AjkVWMlDshloixxkDYj9cZ/mt/flkp6Rs3jftwxOQUG85NXpxvVRzNtzj0RHL
87Ei8uaRoo6Ts8h5Yfb/QxEMzJTpwRSb9X/OUvPuqhtb4NoBfArPzLzhAskpkCMU
P0rzl3Ah0F8Ucvv2HJRK1Hd76vQ9pTlGMqxV3OY4B2U5qcQcW5TZEsRVWefqBNLl
mB6HtA6VRCWOClhEKQr18Zt2j8o5WXnHNz4KLcZsStyNfkq72eKLXetVH7kb9Coh
uddvLANTfdzKgr4k778B3TvB+ZFwaICdYAbzKKmNaAzzDfX+nQI8sv2smB1R36YG
y9ki16fgD0dobFzND5CwMWfF3VoQ8N9EmFvEjrN7L/CRAX74ccIOSsy4BE3SKGG/
Fy7TUyDLKb6omFJDidiUQn7W4uxxQLGkgKdefs/SKFVbLwMse85RnTfRttPGPnWv
ndIzyAgF9Ezz6VHeNiv+KMT11qQClCg92xUuficBc7qH4sYsl2tmIYmqPsC023Ry
oSHAhwYv8SwclWnXFsyHJHE2KK7PMy4TOKsH+cutu4fBo05jVXH08C/zdL7FvCe8
7as/NdYT+vMN2o0rdRDnGWB0AT8B4i/WqDteo8KiN6bQgu3Dp72tZcNskLC7KrOW
LD5hdcIcpWs5tzx4WSTzakuYjeOhJrO4ZLZ6X+pIPTYivGVbDKdfrhXpNhI5vHHk
3itfbx4clr0aaXTeyMSNi+dyUS/2eLzqiLJw7YUjVNvCnOZoC+KYU84S7Rlut8bw
RGwvOqKxVpP0E2zJ/a/gCakwUX3Y4pEBvVOoLWb+TuknmbcCHSFsbpk1RQ/CqZlE
jqeOFi9m7hCnEr3+fV7TvAMphGYnO/j4Xn4Bw7a45DkQZrdBgMflAi8K+xSPWc3Z
HQLa1r3rhYvl7WBFtK8D7qS5Bhu/pMUmN2ocvxG/cbWEnI0eGCvte966rlbrMg6s
s37RZBWxtOy22HoaJ0GOAQfEdEQh9bzU50mCnWFSdyDGutzKlAi9i3CIPtnZ7jfc
WYofeYxhwFwPBAE41md8ZtrPMFWBbkfGYHTavknX+dNw3U2a7+lRiBCkwl8YTrRY
k3C+BWq/AI4kkDucEV07+4/z3ezoBirUHRxIwyJv7p4nKs+7coBM9xxuM1028RXL
OSLYV5xsKJuYCLBSM4yZO+zVklZkMzoJj0H/iEcqfh4babdBMtvntZJR3b99uMNd
lBVOkIpcH2aifyu/ktffpFeQ43LAOrbuh8KWFm0ankUZVP3c6M/bZGgUntunJ/wt
lrTqhweX8ApTzz/jxbtLi4bsKkt7wpqho/bKYL0XpzxKASeh98JXgceGtBvgUD6f
7l//pmXC+TzzZTdYDLurZ+jxjzRpEdspEOEZxQTFeHfIji7XsCSgFvAZMSGsvIn1
JALGGxm+29EWtTsvqMz/kQLezTgzmSfYdKLoQZz8wyWwkAWL7Zxs/aodJZ8uHWqS
iIlYwC4CjazH1rPfCS7LIfkTUnovvi6jlSWfgj15oabMtrhgl0JqWYHgIjyc/VNM
GfPRLLrp96RD+53NTyLlki6gxKO326+1BpOsX38cZOYsR1l4rHmaQlJx7H/0phEv
rFJHg/1vcKEo8hvLJs9XNQtqUAS1v7lMJE/O42fY9wM+phkNsEhOfX2RKa/IgwL7
9I+la5QPLGxB8OCrymtcMVpCqRQCHwEJbjw1Y4+81HkYbxOYFe/W5N9pxq48bkFv
k7PeHc/jkmbJRtLuMJ8Ci85AW2NqRNke6x3XXCk5ouDttmQnuLIMQkQ0N88AUMYh
egWrlbjVkQbdL3ilulebfLBokoC16XwgRDjd/ZlH86q8sDlDyw9JP9j/iBtvMhXO
6PDA/wQCLPlp0NENO634H8Q81S8QUtdvGq/iEgyKdXdoA6k564ju8UD30gLSHNDU
rQA4LN2BVyCIfVHSbZNzt6LcGry54j/bieVhkTQy9IkzXjUf8F8h+iIVTXSinSUB
Oh7Tv3OO91uR3kcVV952YyZDp4ipcik+ERMqUFQWnx5CcBPMnDKc50HkaurVB6EE
z7I/yv+RLGytFqbqLWKZZJOt2x3ENozPbwupeJFklM+VyhBFgpArlC3hQm3pxR/o
48XnCGveYuZJue2vwz7CsdS2rtmSRm25rzGG3TZJXwHyBagLhfuIotTZV7yl2VVX
GLcpv+gnGE252dEu5xhXPqpA9cAGDyMluNuzB4myPMJaP9bRgdFBt2DpjFSg9twf
pQ5I/bNzTLdO0kgGj1rAA2aNYXTCYK1q9V8VAnsnMnljE2QPdTkyF5z7bSURf+Dl
U5Y92iBHYIin+QmsMoHMcsHwTGir9NLLUDUs4D5DHcm1upPYPokm0DqZukbv8ULK
8WxLiFu1/hl33bHfr640gYQWkmkab6ZIIeELC5jT42zGa977u5hOTUuQOayRWhWO
fyDs9BTZwuZD6pyqaJSdBDlyQ+0RtiqDwAHYkHd/jjEy2mW/0a02sIoC9aBbA148
1P7MubeUlXcwj7XQsoTYKwIoX5th7tnIumrEgatTjUR6GrONLj8UNbu0ptEhiung
rDlHeKgbwgIou/jsBZ8swGxw0ZC0LZW+jp0P1iDwmu//tDPjqvZhKmjCYaIHSm+d
fhr6I56nmRT1hilR1jGZECCuWnwteHlJ5kkixwIW4qbS1JPmVepAgh9cfPpZsJLF
nyZxX6jvd7Xa41ifJgOeX1anP22tzjbfjR8pzPPXOnNhi8+QL+COLLHcCSugCOUU
qq5lPrIua7IujgxuA916ZHhITFo269WDMisLZE44qYeh+RBvZ2sI96Mr16A+kPM5
QVgehWL/b0Oz82lDajzwGyNdVNL+/3H6vOPnesSvtMxBvUnjcgyUcepoV018D1C5
rdjHVC1rU/hfKtHYEjybdzj+JagaYfD/PWvD5jURcBpzeZmvq58dZ346Ms8qPzqB
qYTgFcIVcgMFt8PIV314JI8y0Bmdp+q/s3Y6IaJ+Thigx7MYjqXHYJJaQUGp7UJx
e12RMBfFdxO2zK9RGi7rhyQlz8CTAXTGMNba9f0v9nCqIvuyzerdKwZuZhIjjXgn
zswdsWRAzasH+ClBWbR9cPxl0Y1Cd4c3DpwhyQRl1HqKn77m+tJjTaLuGxDOksBZ
6kGJgqJK47c6X/WiBM4OwvAVl3GdQBrQ9SChKew5xG6tUXXvrnjVq+CNHARJiC44
JyeICOKrWKJ9LI2a1hOLq9cdcZrblcXmCgXUdu3Baqo2kx93fg+aKjXAPb4NPzOJ
SBUOmr74uaBcDJgRmSrzyeGM17UqhPGNO91H1/oavu4wW0nhh2xHR4gwFgmvfL/o
VcFP89DNIcLVXEH2fUK7M2AqLpD2QHjcnogyQ77SesAehoeqNIwCjvNXb1/ILkLq
V+oUD/NNOadXMSebjDKhZ7vrS9ZOs0t0bL63yfXLkcwp/bNNWMlvEM6FFlz5OTEZ
YrHpddhBwBGSgytRsLnnANAhMsPtVpPTlzFcPhF4X4dH6diMItN0q5oxr0vofdGE
Gb4z4ZV96BqAiPC+O2Kw5Z+mZ+bK4T8mlSttPHJxtRmYjxTxM7wXQncNzvSdZv87
7kIgp9B/M8I1JJBV9RV3o+enlit81JAn6eRQbSeLjkJ/cxU9G0MAu/kBdWcfToXz
j0409FJ1Hi4rx65xzoxollAkhyN94vtTorJXCVaJhMNoey5iUbmnAIkWj/2qFVcA
vsfz/QIdx06OBCkXGs8oqKkkg+djKMxJDz0PigDz3Mg6pYkCyWlNxX+g9HNaYYdv
CLc3DDA1NnLMv+vBA0lbrT9ie+UsulJ7E7610EfjaNKWmX6pqJbq8b+ASUOU8WP0
Vl6bMq0QwQWBoZwqug/yMpCm+VYlDPvNFpNuJqHaWnfkNjT5Vce1nuyxTmJZc/3F
197I3wcYDU++L1K+y3eRoEqpGU22B3WQbWheBF/Ifb5j5gDJp4fI+TCSwGkOopSb
2qUn3EGjWm4zIpmNPeG7PEUNDpu3plsUgTqRk3aiWOykXiUnXnEc/DVccPJoNp6K
NV3T8ofbLKXzT3TvpqmDZ7CsXjUXPX7DPAlw2NU9Otx3xqtuIsGEq4x++kTeDanv
x8AoRe8UYWzRkwkKpIF50tPWsaXwYvuuDeZm4cLIm0qF92cseciuzAlk1TfbCBut
vrqH9jN3TJHj6mjxDG4TagdJO1AjPMB3fOFblV/blwN6Nzl/Y3dAPVv4dc+852t1
DEOEdTXR39mF9YhJE5UuB3U95OeGuQsMSvwXne4BTySF2/EM3r1cQvNFLEf/rAhX
zzngIOh2UEYFw38jMQa5gPDis4itUxZAf8KhrePrwnkATYG1gOORV9yqnoC6bPou
jUYvuGihCCZ0Q6WXJ6fOBaCoZF03MMr2UN1dRwuWuiHHbDk83lFYBNv5uMHUt4UR
rsFJmzmf//Gwa7GvrcKG0VK7BBzg+jaV24oEUrKnrpXcCd2Os2/iUrv7ep1WfXQS
2PiD8Ccax3XoPGeNE9aqmwVBp88f9Y8XTw9TWp2qI1wdkNPEuT9ggMFTs0HfobFm
S7+6G+JN1ppEx9m96ibY0F6OIBigp74yLYUzActGS4V7lhQ40+mHJTbfkJFMNoO+
HS22vI2UtPY0WqdDfewtuTk20y6ZO2HYWm+HSRjZwszF5+dLVnrU/Wawjs1Gw1Bi
EXUtAM8ER97i17b7e9HfY9WpWuChHFrZio079lAr8esIhc7b/VGV+ChfNc9JL5iN
/I/nVGEZ2DOi0eBzItBHXC6WrjuagRIPBnuAzIRtA1EFEqxAehwruzUDJzvCqNFp
QDBe6Y4mFMadQrJzW2QHiPUTUVrAtVovwHeWdVmWLHfT9hHqoCcvzmDBbZ3GjXGH
7/usF5H1Gx5o2D8aaGoqWB/XqH633jymojiLmFc/+fa71MFiFIyreE11QfAOMrak
+kUtkgxqyEK9f+isgpK64q8c8OKXqY8ETcpFkldom4WXrgRfOQihb394I9kAxg6M
awx7sK+4SMyqrMJ9KJSpWoP5iEfyu85LVJ/bucU5bpy51lGw0JrJIPZEu4iPvZ89
hL4anJd7xoq4Pvrg0C/LNbPv/Vb7KHzQ9GniuPigXJW1gxqt2WwOcgkLvB1lLfm/
Y+YY64PlCVc5/vUYfE2SYikYf6w/+L6vbm20qB0cMbVeQhSoCv7Pepfn3YW3Sjcb
SzJq0igu2M88BdzXlIrC7dyCFf0TWmkRWdhjCucdDODcwjsfDjqXFVKoPzEqe4Ul
FpN9IjFLh8ER3QFnLf1V9WNLuHf+bjpgX3AdqMO/7bFyQ/rhyP5h41GTW1HBiaSu
Qw0OV+b9KMsxdqfbc9AAl3bGKuaP8qKBdDhy8MvAm2H2d4dgXIq8XEA0kuU17X4y
WVCF8AB1Vte1Po+7uQiEWUHY3cjaDqkhtGABUHAkyF8F07J8owXZzofEZ7B1yaJR
S78q/xb9CWM93tessFCxHqF+wMraAVyx8FavjUnkt3wxWDahjSwdfe5VpqyW8TH1
mZiAIlH1Pgn1aHh6v21QmB2ri+xLcND0XrEf0Krk3H/mL0RF6qN0yHpz0zXcegHL
xtrz+PHSB7FPTSEdx7nMK9EZ6e6z3ADt/7cdXyxnwAnS4+E5kzAPrmrmQPYmdFEm
4zq8Ikxqi+kmUiz1WNVWCB8bA1r4Ci/+Lc9wM9ZD4u5McUzJjEQxfjYOuNpATeVj
XnO+eah6PAjoc+UDuxbY+VvikOCq5m9ZnwamuEvy6AiFXwin9qPr6ltwIag5O4Wu
SljJPJ9i4kdZdj4MgjTXkPeC8ntHEiqQ//uqkdEL7N72ZSVYB4XmnfJbNL/LAHsz
c1dGfUOiseBxbvpfGI/TxX0tMhQercDT4+GsrOv8tfEjvY6oMUpypMFQ9kTarbwe
SV1VmtB+6A4Nic0BKzIpY5K45jazY+5pFm6GA8vTM/bdTn9QZ9PuXQ3mwZOgrUON
qsuMeFymv0rT1n/QQfxToXb14mpT/Aw6XYw1AdiNtr7pJK6xowQDVh5ba9szyrq4
exobMYuS7sMw1YfFk2eMoiXD7B6VsWw0N3jD3BlAV1wby+z63okAbYqHK2FHoYWo
QOUWXaCDWuUEnD9pC949JxzZac5sWBcRRKO7cNt44vaX7QtE51KFanUv3qvfPG4w
DLx39U4KwRWfZeGMM+cNES1XyAMKb6GTOawZpjEc8fL02a1mZtM/QiY5S2Pfm8DX
Ly7tvg3/vilLGFjZ9aQFiw4MhGG9IM2ikD87aOxSikAF7kW3ZeMILisNjcMhm5Tz
xzX9OSvoIXwKY1dZ2qRSHVjIWErlZG4pjXpttNNE/QSWXlpL0fA/idYuqAXPHiOt
mF1xxDK49GKS++AfLd428hEmABtO10FhMCE1/O/1h7XgDidQFU+OHUOefnZ4xtII
255YgTeOG5KWY1ugu6RMN+/nm+6VIk8JE3L9A3Guus/IO0EKvCnIIlwXVX+i6GXu
jVJO/GlEQ00Qgl5GCCnHX1RmC9Jcl7zZsoE5FwFz0IEZ+aJJGmSkQSGLGt13fKld
gwyfozIPFidWkeU/SLqpfqHs4QqlgY/7Y2oBjHs+OvNSlma/r5yXqXgNfSUHnMd2
n2WwG7LhwGiX/gcXpA6cRUgOmi/rIM92Xp1mm8WZG0HQ+iEfSQO14uuG4yuNhZF+
/hXo6k58AL6Ri/0nLrbi15Kkj3z+kIR1+SYAyoh0GIT6DdBJNjFQZE820rbq2VfY
8y4efi0NkUJjHxz6yqz7vny9/PN62aRo33GjGd82TSsrVNhq+zNuEYVUC/pARcAv
LuxbHhpdewd/IHJFQ7upQqIqGAVOW2tSNomeWmW7e2Q0Qaj3O1f1NDwkV7eJUddW
DQrnCBioHqwP+aWRGaEYO7S+U9EM1KU+yTnt9cES0jLohyZkiNBzcdDuE/fMAtxP
gitkY1S6dOz8jLugmQpaTa/CwfJE3AGMcy4hhVTZKOlhgcTZ/LEQzFie9jcur/Ih
pXjbHT7irxHgodOmO1eNG1X+KG1YBQgTDlEUkDcqEnKi5leNpXn6m6fFjrApmTpy
NIsdoRxyH0Jm7y5ocHPAYacNTPfTQeVKVkUBzrgxIW+jLgtaQED/GZwo9lYEhG8B
tet3oN/KqBvQOSpxHt4HmP7r2xNqwz1jcg7uxRffjZe0EgTZYk3Ly0Q9Z7VLmn5/
f4Dl6CFhmmqxAtns8gZLk7e8m5ddAJ+XJgTl/2Rx2t4GaNbr1M+A/l8l2gIBe6BO
nOwfX+VwiQtLkOAvwJMSnxh2X4KHG9eDs8+1Uyd9+ZrT7PY17raXFg60QU1F0KJh
bYxHbj1vt3CPZasYpMs31q9dPCxk78GuuDAXmUxRLV/WG7oJDt/HO2NpIsw5TJjS
WOdn/G8OyK4DLzV30KWWxc43dg8ARbuwk4Djb5MdAmbFRcvsbrrUdKYPyjDDSizB
1VfSxZRq8aalwMogpdJh1meyNBBNr3WSPl5WtNtBjamqcxBrULxhqpC9PW6d99gj
MQikISAqGLmlE3mtj9CYklqsmYpW9dwQxKE67BW3QfyAoBSvWz+Ay81KXrgkGZbq
gKuEgFmbNNZI6ls6xdI3+6LkvmBW6/VTAQdPMVhBdwfQ/S0cwH3qJwuy0/HR27P8
W5KDWqwZogMBlUzS7SIBfXZiY/hcYVQ+FEDWCKNQ+Arkj+OyWKJr36L3WsgM/tep
ts1Yf5BqS+i5HGGhUXg6kQzESU1AeqR14poYyvWmgIgKTOhfIiO2WmadW/Qz3mdV
4ARyblSIMZ2AaMQ/a82sbUDPGwK6+3hXVXZdGWicN9fpH2h21wu7mQ+icrexN6XP
xzmm7WijCIrsSlcvGQ7nFVeGWJ+u6kbkI57Ntt3pgLTxAgcC2XvpziOTHz5ZFLdj
Ixq1yVn54HU3ZBOcGncJxpSxPnLH9WJpSYfDYDs4+L8tn2LSiwmu5RnLV6V/qVVK
3iIBH7Z6L3b+fDZWsVUFoS6bLoLjDjNfd+SqJy5E7hKIYzqNnflCxj7ahh8x+3DW
4Pw8eDzlB0nKb39X2nfg3qj8zeYwCv31GJd98YK9j3WGNeh3StohxhCjX/V/oBvh
KD8UwFjbC28Txn5eof5nyefhFXthFtWqRElK75c/bZPqXTdqNfOCV8BsvEsNyV3Y
mopNBYuX6g8sVMYDgMW09sxlpUJG66FhCGWpp83zQMy5A4DPXylRrLS1O1cvfqG6
5jcd63VMTQq1QrZdJVGY0U10elzdo27a5IsQnPaK3MRSKCbtM6Bmws1Tz2El1pjT
2K8DDbxGz0MoUM7xpNSPEOG7+taUwN2zG/8CbVVtU492VOAs7wCPBdINopJ3Ct8Z
MbKBc3b3CTUaksIeO3B1KNXabCSmDfiMQUrqD2LYHuPRfFTBRtIVpBfnXX3XSneW
SrS3I8leTpjeTMvNSqCFxF/B+4sLMf/aJ8WCBdfNJkEusZutjuMwysF31U0zZECR
YkeNq3B869zUadxi7FCSYvy5zMBtuhM9Yw9ELcjuTzAhH4MbE6xdb1cJ/jrKpsvo
gnhsAQROjuf5lfSikfVdhTPtyFvL1G1+CSAWNNAEmDQ93WOdXnyRGAyvNQpnjpIF
DYGPBkJaryXVn7Sv8YxvM3ZOAqSeqsyyfMP7xr2nK1cerHYnNSuK3oJSKJBWxZAR
0/Wtprbf0yTywVxHj+VMgqiS8GondoXtehe9HQ6bdzWRRD/CqW2j2XWyjwT1idVd
H4AGlFhbubtS01JUIpiizCrv9TzmbBf+uyAAILKkQdpRWoIb/hH0+B49nLu7ZeMH
8vkTSPdg0YfbA5xX3EsMb7gciKQn7Git/VLzaYRRxHVTLVzuy+wuxX9M+rDF0DCH
1juw/vzaWmN4ECuaKz0rJY6geK0J/EyUSVuNb8bjPQ/qsnGe/0av9NPVN2KNYuy+
ORlJYYNCD4i26AGX1t5kJWnxgLCmAzJlBDAxAJHFAkyZ7HmwQhxCYwEl28WMAvkS
4XvBgCC7wy6K/TnnDEMuLl0MDy7FGcs1kgImS+MW4eHIw/37vCC5S4Bu23JEKgfs
w9YTpWm2/0ggPBTLugXdbfs8ZdgdxJavzcvjFZmadllBzt+3BzR26rCqjcj7dO5h
kXRhlbh5WrbWnbnx3rwXDl3yCSgMbVg8jUmpPvTUHlUtxKfb5Nk2z+wYOw+RA6xM
jPRv9c5XcDCHdvIRt+bnkEPyurgO/IsP0qXKhCIxitQiihxNPBApMhMj2eE6/C3V
igJJbd1X9GVKP8L0b67yzUeSNQASCYjqs9KauQ81zni9Ozsb8SCqIKQr0ycJ/9s1
rTk36EPLbpdjrxTeNBgCgfn4NSnQZsuvAYkW6BltRslvG05sNDu2izRGW3ul20yn
dDQOmX/cMkVc1K6FvGdF5VEh26Np7abaaFST4BZtJEYtYLmd9SNA+fl47E/uG5rK
IISzE5WFAmOzPptdmv0v0yNi0MGxlWwkUDWZ2MX6PIJPP0wwmU0Lqcz6YqqXrEzi
nOf0RJ20L49SJvFA1nH9rH4+Mrmq7GvUY3ddRwDYnL/8j0G9DhZU8k4aMWT/JOT9
EgUVu+YTJ5R0lYN6HBdOshH7UZenAd9kxsqZixwS0Bs9pP/QLNbycwevmU4raZCw
NirtpBPF8nJzg8oPyctae7Yx1lgDjpoCd2C759d6e2WzlM0Rd2bN1RBLzSZ12bKf
kvVmDp6CfW10oAWaz9GFqIWU6XTE9/UnZE9sAo5LsGw0N9qYZoXSJGajmjMJpv//
o7w0sEqvdGIlufl9wrJl1S5m0mNnLezJX79axLfQjfaE2x6elRKt2IAAJjq/pYUf
bQN4usC68GTV4h48FsI27Cm4NPSji6EXl/WJMJnSX+ykpM1YoH9izOTQ+miujhJc
YvZsCs2OtNTNIb9pjHN+HFRLVdq4Qt4Zbus2KeYAVt3LbVpgJ579pXWPfJu97sZ9
j9MKc+0TaqNcopKgx2t51KZ65jzJMot5dgy22gIarRz1VrkZgcNOOJIZDEVtgvmf
DtMJBPx1JhD2J+uEsIsUw9X+4DbbzWg5gmtCvrEqSqx/tbMYce5oUqHkodKQSHTF
A1SrlbvkjN1L4Yatw1bCMJwNNTjslJz39VTC7hgeks3hHWesCYD+GRtsrhIBXCaW
iZKI6+7Mnedfqe0KLfUGzMmH58+74phZLodcPRkvj6CrWXHnvGuY8bzAt3JQUggx
Xe7/2htHWPB2qJxpum95MhEVQjLZO+v22OqUoK535GCSBrHZoNczWIN3M2/Lgnct
WF5tJIl3I6xdxwUm2ARL4wkR6fveDOYRYSHIBmvTy/Q5xYQt/iI1MEkJPRj7vnWE
0kSjg4nt87KFCY3V5Ry5fEH3dfGOWscITvPHOfrVyygpM6D/VJq4kzDR6XpoweYg
ABAdQlaPKkn3Xy0RTxMNgxf2aLQfTq1+dkU1jT8KmYDHbvnDLH/f0kRSTIWkMqP5
TNC8FxHaCWZ862RbeXOLa790zowNi2+Cadp+gam7qf9K4GUwLNea86+BGux/jobo
3IIlQtqGyF1R0YxAqxy9BfsJEbT+BvWUCZL0zg2ELSzqKjJF+GAmd+lMFYwizaqQ
H4/O+DAAdPzgWxpcoysAqHzuiNITAlYmefNCCncsYDi/wDLw1D0y+ZzD8CkYcW6A
FHn0o16UMj7eTLT+1qaPOFtiaJdSO4dL1Oy5CgM8F7QU6+GetAHlNOYWd7qzk4Q+
hxOg90KlNPnI1lB1CVdtAdT6le6N+GexBFm6sKtrjW413P6Z7a79ryxV0XgwDO88
jIhYVjHQ5dfikG20eBZfBslt5jjfWknoWOPl9eQgcbedveJynYBohX/JgFHLoV4o
`pragma protect end_protected
