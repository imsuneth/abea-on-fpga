// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:58 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fTZw0Lw3zFonRTRqTaHr+SpMvFfDehK9aXH4AZLZ5gvGo2jdleyNnxiA3tdJeLR6
8yL7PoPxJLE9cTTaa82YnxSDc9aDEatzcb/OnIc5gKOeRnUOhlxPNL1MuaAUrcnN
cGCfSlfFThR9yhKljR2cMNhJkv9t+5AciIquaBq6k58=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11648)
or5Bu9NcgDHShbzgzAFBqs404RgFPZ+kY9vJMjTuJo2iW//cdhTyQlCDujaNiJvh
CCIT1JGzTSjVRgAWZXluKF9ClN/P9dD1HMZmWZRXwfH553lcAVdjx6HLyI+XsP+H
x/2pubn5SVz8pvtCSiNgXqlnOiWtaBxu+adicNxKnIOIm9WqeWzF6ccUQTIDL83l
gEyevpOUniZ9nlbaTt0bF1xUapJCUtuiZV2IIuH/td8PoRnC4N1BGswQ9KBGHa/I
kxe6liwbFAowRpCx+03gdvOfALrYoGU15cD506TjMM4Wj7bcU5B67gW2G5evkCWw
+LNArq+RAPduRA793m58jMLopYQGByenzdAyRpQeizI/owGxuAMdcWoBXJFUkXqR
FpjGG9mqJb4S9hgzRwsX4/GlkHI+N7PKm244ODfMdgnDftYkd4COwLzGdoa1FIdU
u/tVVnJzG8KK5OAAwsfv5+d9YpSYLTiWokRPCRULeQ6sUwpATSghC3lWmao6HV25
5i3D8VQ2rasb2wkLPABajyMwv/Rq6r0BMGaS7ZuXsSnYZ4ISAECKcbIvqIe+9RDH
mfoAsNesgLGKYucIJPfGCsuCc4cjaucCH8s76gyR4ynj3tAAlzpIWWP7kghKBaIw
a2mq7di8P21AMDDoXPDg7DjeFmBDbTBGZ16RciR7CJ5FnjzNUPuUd3rAyZ0Al5T1
Rvj+oYBKsUIYCo0YfJG2LPk6nuONIf+ljdootko2sVPwUWBq0crEz3PfL94wln9T
F8ka4JudDFUKtDLUvJ7gGKitGzDjryP2PxbioJayT4Le84AGd2whfXN49h0jyEYP
qoFJXTcyZDK2EXou9gTabSymPmidN6HWSAsFdx6D6EtZUV6Ji0Gwl6YX9bnDaq3z
vCrZNmnAvIKPdNv/0vPSsdz1i2SA1fPRDm1O8woc8nFYm320x3qEUWO87UgIYKua
mqqhG5V9jSZ7wuRn/RuRoUHnCufz7dVnlEE/C5Apeskn45UB+TjYYUzDRWDQOu6C
1yddHkZkWd8y79f2zA4QjQoSMPo8sa7lO9lrs1R6Eh3W5VMKNnAvPY4HCpG5qesT
GyxjODMoIRQQKvA01KiwAz8jTs+32n6UPOCwlcy44RM+jLptUQGhwXyMXzIvv58t
397dsoLnDarYZKApi+fxd71HmgscXVhXp1URVSnWoHZpl68LdxP7ecMNKwuPTw0O
5xMCyZYLSyB0ko2pTl8tpyxzPO4e0iOfqyCRTonr4A7JhZiwB/94U/2IwA5kYfRH
dPmYv9QLogpz5oKPQTkhzMjeCbLiDFFu3P635lWvPAaS+nxib311opJwDq8EMT7j
4godA8Zr5A0T2NnslW4MpY7RkuRQbHMqWGUJRi2LSeRbNKkVMnAX0TGO8/xcAilM
nS1zavZvcr3XWLhIy51NurnkgB04JXbKCKHaH6EJRN4k6x9UtqFXXotdx3PjgL96
NEJU4a7aOXVt7m1OG+Zf7bPao9vchjn3N/2G/3opyfweZXE+WZP+OwQuHKMxOmMx
1FRTSo1SRrV8TX1IjV7SVeDYP9sFjppLhdn6v1+TXyfFJULYmoqS3NcSPu1BWaFe
M1hHXiWuWLxIdDQuCahjEDjmxhkE03vtm+iDmmGMQ13uqIE5nX8WIg2GhlN3MWN+
RXUGehRh7X1TJVqHxmo1CZqRNRIvw3OQoxM8oPaaQpsVB+3eovp6XF0wSq4guUfH
hqxC4W2vI5ybsv86L6KLpFxd40oGtq6/caz2gh3qrf9CiSNbhdJvfTllZom0PSUi
U+Lba5I3PYUdWGkIh7aJUHSCXUpriO5goUd92hUU0v3vmxdpTj6dvag18ximqNmF
Rdn9Qz8HmUy+8rdYbLjJgpxX7wmPYIO1fnIcOpTxHttWbaQm3hFERa4O/0+yVLXG
7gyWtSrhfT0nJ7rk65cQiA/9/FXxbG3I65+Pzc7dsctiC66n/0e1Y/qaedO2XtE4
6TrYBNlENmZGq4wnnFJwvpcgPbsuht1WcaIcA62mhssta2HAK2qgXJRLHZUWkND0
9WZodeorykcbLBAYglydwRS3lHKfmiVASH5oskseJh02lhO6aoDHRNnwMsRioX82
Fs/tC2jV95K7GMa2Ay8hjzoYsSDWJOr7msRjP3G/VyN8OIfoVJM0DfPfX2zyTAuU
6ZkTI5N4LMXcrTgNg9QYXy/r+O8f9L/ShfWk6SwSewhpOcjk8lxkydbTnGAqBZZ2
Occd+Of4ba/JKnDYb4PrbWaXrcV705AhAx5S5EfYIaBnRIEO7pNHcCVKI1NTnULx
AwCJXtg/DwiKHD65GI8aFO/jea26HdcRoH8JhLxx4gMtR1wMIb9CQo4kbNJ/dIm0
cbFwC7NtM3Bo2CBnldLvbKF86iYbifTPqNMmCvxIsBy2j/Am4s9jXjTuR3BSiWqh
yQuxDH9vmGVBlq8fGmQyffs7K5GUegYEmsUVuaSkt+RXnVTWgAG54/YwE7gUVidK
t4BVqAI8QmC0pVFdFxCRCz1bxir2WRMwhTtNK+namoHC0IMuwDDeczyqh0bT+i/J
zoTehCbPjX0lhLztla1hjtW/evCWPZSlnpk7hci6uxNuLJbHnPv68PeUtTB4gVDs
9XzJ6/0r9cYBVffM2IghIHg81LOzK0zKcgt99IqxYpN114w54jG+hahfuEh8W580
EkTZ3K91yMV0WdASwbLJgoC18l6etuTgCAnmA6teep2zkUPC2t8it+ODc8RNhMMz
teTa06RBN036Jjwh78T0JFnq45aNj9q6DcvzFxs6x1UhxzSR304Ap1VZVictfzBz
SizGZfYk5Un7PAj1D5pFYhe/GpAqdcFn72BddcrWwd8a/8rh+NWGi7JwuVtFTnji
MUzNR+2bKahelPMugg1TDXdSyX3zsBRB3uw8+wxzH5WNVisrzWNKFt8WaAd2IV1O
vCfKs3qaMzqMEaMbKCHZGrHO5rdxjKn8bFdubAIKw8RYjJvwnK99laIxdcG6fXTk
9ZwKiC76BFjto2Tzt2VAW0ETp/sPWT2mLbNA7nW5GOswDW6GOWNRr3M8qw4MROC3
96c0trnJJcREwGfaUbPVxWm1lJik2ZgeAA6mxlWLGJ+80Yv8dDGM+kTd2h1QXMKe
7m36yYnUhLm+xKnvcA9IKRokSeWwM6iGSBfXtZ741/m8NNsV1IcCG7wsX6hwaDJl
vX8afZRyPrrcwYYnONRooOfW30hYu+0RAWUQ97Efn1xWZFiT7k3HUKkOkXkeDCZo
EB4QmMLZEbKzwCHnqjK3xG7EULS0vcKHFkB0A+CJrFgFIUg/Q0FBQ9f7jM9bMywz
BcfhJnA2sLETQxpzjcVWGHnp3+M2Fr2kQ9fthxQfMus6dNKgQ4s1VzDlP7AK0hYX
Utw6VfDUzeVHtlZ79ZJ/VllfawWy4OC2HjsXvCao226PVg9hWrAl7rDqrorZbSh3
C/rfbdjHNEgGv7AsKqVYsAX2+dfvdkTkaAcmEw8Ze0bfJ657E1cYr/mq9gh78DZW
faRzOUTujOBcXKnij4B6ycv617bKmbh7jrxxpbKsFtJOF1ZZ9qesAy8ad1smYkZl
hA/N8uaOTR/TDhf2RsHGarooINM3jrThS5AsgjOxh1o+XH/VLXgQH5FB7eoOdeb+
2d8jB10SwyQAW3VwmowZNjuJWmyf0ovRbO5D627TYyGJaOCg9mQYDYrXhyJnwbA0
HvHNL6L4IMh9OE94FK6pEcrxSE7gAGOAsU+pHeYmj9W8mzaIzhbdoos1oVCki414
+17WwZGsy87Arl7In6hytDiSWHNfprktFIhF9NX010LDV6mOFJfL8z1Oc4/82ZAv
kLFY8cNxrGWG6x88lzrTFvN1zCNhKgGLPazjp8oYZSxHs6Z0+Jnk4JYmuWIWxp3J
t1zhcVCdUUNFirKIKtRLKNzoqFvXTTlbeoRcfhHZ4PHR4b569jxmbvMxg+hVylR7
aQ/FzOp9kQ+tcpm2G9CZvmciKoNXUys2CcEWSpE9b9aOgPIY7CXEBK7ZUde/iB4J
Z5qs2YmbABVnfgamAgtoL+fmZoV6AWfln5F10S0s5xPLlioQ8eXt9+R0OzJ3DprU
Ufz2Ycr/Cdlch1P1Ot9p4d4wZ6KvtOSOf/+OGYQfDPbnCGOJyvygKfYDhTLmxia8
7hQ+AoFb/q766unOLaexnlRjkdu0TAgGHRU9mvHDgDwLTU1lnizwzmpBgGV2jCSu
4sER9Ry9QGheGHIpVjY1YoinBbKzAI4JJiQxtZF6Sg1cxMbVQ6ROP9Mzs8mLL++m
99QzX7cyq8xeSnAfrWgZXSCqYW1ExAlasPCIa3d6zmDtEJXfMCQWW7bSSBa9bJSR
6Ja2y/iZPcTiN6EyE1ccD1yUXnBbAZMb5RdnQj0hEM0LIfMst1vySZdvFZl2D38r
0ZbQdX83exG0gYAQw01eH/D0OGEkxKkBL7xrcQJz4IrbWRCVn08Yr8lycIYBcIUG
zyLQs6iIOqPH5Rw8VvKe+lHuKd55oPppb2DURCQqmEGLVdA21cUsw+fI/blTWXd9
NI02Z3DD2ko/X56/jxQKors9uemnrHe57CgoheG5OZYLgC//X3CgiVakRjd77h5I
GMQ7fN8FOnel/GzvgElCS7x0BtZMucY3V9fSVzOrTxdNOQ+6NAbfSL70C3PVf5gz
+sQNeR4L9VGfv5aui8YDnW+Z2dsAjdNYHro7kUGo0UEozuiPt9jt5cO1vptMm3AR
lHQwVg5Jaxq0VPGFpGsCL0MjEN7EhyerKei4XvUEBojPunWCneV6dJIgNwoHwg/s
HSkJSJk2QL7EzoG9VESkX6z16P8tG88nP/vN82Xc619NDxQ0oUCyFnKQ9CbxFFfE
nkphhgtBUZutFGm9F6/SsoXUuRJJ6YM1KUfMsSLYj7QaxiHUWc+G18JGwbBZL9Pk
GVVFgBaV4KodXmlW6xLngZn6w531wiRK7HE7fH+3xZJ7MrWncnxflLagt4kXwxmO
hj2f3r0ctz6LZD5q9Z0lHfkOem76BTOW45YBuZp/MhjyynSxhvtkgkw6u0DxihZc
Uky1+QxRnGAAXM1fvDGk07huEYjfQRZZjFwdHmh+dvhwlRG2Wp4E6xOtvw05/6jF
tvuOhbKolBao/1Fp3Ba4DwwfuiDkBo7kT670qcmcn+LYglpDtbIp+j0Y8MhU8+Wr
p36pUL8MiPr4vBOn3Z74X4YoNbRqGDgCxcso42EHoRmjvUuHUtq+DOwmiVwx79Os
n/VTqjpdyNrTSbBuZoezQ5iM0MTwn3A3sLGvtubdT9ZSiWyr/T9DkmcC+HXwhIxK
64Dcg4QfMQUgPsV9rZg4fCDOcd9dkOObmcTcoZozTr2DJV6SSA+3vTY1I4dgdJcL
qkt8sCR0z0x1XyFaGvm964rUILcxHHv2luW4zTRNoPLDuiGfDVaT97am3xbjh/on
7hPvtUx42az8JQoSg9SuK4MQk/2j6IvUVQ8baKcKQa4DKNu5hnddN6ml6pMdbU1l
D6n+Gpxdd4P+9WzhKCuOLxNfAjXIXVl+KSWWBnFOUR5YMGDMX5wy2+yjmeH2otnr
yPW/wW3hnUGth6J3wIOxP81gUKCXUIXXLpxNX2n+kC42rBJV82ZpucvdgGE8BwN4
tHUZ7zbRlZlEVhidE72vBhecXp2zjVSV8zJq+lzM+JKyr5jBFY5B/jm5lO7vq5Zi
xQ6Uqs+3F5ind9kXOTT4URpcxdMqK7s4N9vBo+zWK4uriX9mxshBejB8Wq9BauQ4
fcgxASlA53O7DoKiA1UjQiHfi1rSBIRFT7sq1l9ZXwGvEo5iuDPEu/dvRrTpG2M3
KPUJBm47rKwwQKymN4guPUpGqYuklPZL+44jh2aWBZqsSc68IZ3v80YSlgmlJD3m
04iAqs24CVvD/cW49qrKL/uNuJdejjNATUAZ9oTybGoIm4yxt8FW8sc7GU4tTMRE
nex9gLunp7a9GV5gTyzyRguNvDUOwxvdxRYq8cIem7hlwl9Mc40ENNnVOnRhb6J0
nFmjWRAblsUmiQbqZVkDg2Ze9HniQAx533uOfS+y2n2mdywS+mSKGXPUqm28faIE
a0YpGLmhi19fkEFJeHUITBQph7Mn0iuVNczxRsxRsM6hBA7xl9ucuk54fShLuLuT
E7GnBAOTJqz9vqCOoQz9EoCLuXEPEF7gMWFP89hRsUzrc7bo2P+vo0i65/KfzoLO
jzJf+SjQIQdHY3pxnWdqMsEoHd8Hfyf8cxZjkHoFhTFOrv9aciQvqNdZG08B73yx
P/xpF/uBmJvZjGDGATMKI3xHvCSeMOi82a8oc2LGTKjb973T0h64ZcuHRR/It+83
f8j1TVVnpkE7HVhgYyUyMrOvmTPGp0PxcEjgH8xJOSpMeGeCykkfy9zqH46dynxX
qI84tIL/uhNKuZ9qkwoGe09UCgCGY9xpLwvhynW37Fo8DcNySdf2DSBMRiSJv5Is
uwQOvFOWm0zW4c2tGoEyq3gnnZkaj8oKO38BHn1rRhUDsu7XMzGYUj9olpS3296+
g3TlLXaoDCmiOPPkb3b02ZiQH4LECOoRSyZa6HN6Eufxo+d3Mo6xnLYrQxH+vfvR
FApU8SmcBq54Kk0zXyuQXVSxGhbp60GfLolOeiuN7v9QA+ycO5gBZeEJPmtZDzER
1dWbUNNxCV9yuQVs/B6age3vA+4iCm5nIcOQnPKf6Q7uN7jTOIjSVwBmWDPwsj/K
D0L0HW+rSNMKtAVdBOiYBCipSjirslWPzZ/RvSxCNQko2hSdnP5s9jCdQJdQE09N
mCYkJw24CXHmQfhS2A6imua0MX7GxglkJd99avHmtMezW0Wk4KPKfwMyTThV9bLY
s5k6SGgPldWpM1pxzBZRBzOICpjoWCv9u0WIQACUzr2KtIn+NN3gKeXgKyZx3NiF
YLuT+SwWnzzNT7Ntb2kmhUZBbbKc3zydDUQoN3F2yNpeXuBMs+o7QdpEmUuPAfQV
pvicLsuZyvYco07D9DHcCY7C1KPKMCktfuAWYktZo6mcFBOzqTT4djzsXga8ASzO
HX6FRD7YAdOVHzeecKV5YFsY6R1rG+j/WZ9CKQVWg7Ix6vUzkI6wddLwMBO9gsqj
gGnrWe6HLByoWLsi6p+MrinVoUu9sqQpz5lEdS9cvByq9R1U3Kw5FtTAv0t9nxyp
t4McSJr1ICxh8DKJy6upPx+2darEhI4/ylN+yi8LM9RcctGUI7wdYdMr0ug1gdlw
pZRAq4WqOcimbVMMnYptf/uOUGQxQKzWtdIRfpX7Lzd2FZkDlf51nX0D6/ylJcOZ
o1KYJQ9zZcH1+WJURmy14Rg3EpGob78KzIJvHAyeGCZylfRnPDTOUIGPNj1Vp9Kw
UyEEBfC5NKWXzBHFrm6cSycotPbRHjtIB8og1soDQ1Ahe5P6l9NLKFrSwuZQMKxN
JB+QIf20vHTcQg8o9h5nSIFCbZeO98Qm3f9rLtPKvYrRhOhQBVJon9mmApvKaCrO
U6Las6PoDIHjUJAd5vPYP1qKOMcX77+WonYNQK53TgTSRxX54Z1JI9O0K7Q3JHOZ
siVsoBoDGoZo8rRoVjoNFXOd0qBkYtH4j3vQvpiOgVn0qbCL3ANAo6xdB6op+oyt
Kcmy3aazhsiB1I90tjLVG5PoITjA/7c+W6XBJU/VqSavhQW9M1LgEWc8MTHJnkS2
99ph04sJDrBj3dir30sajxOmDcJFNN4P4DWWT93yD1nhIPLApDLfomnoWnKYcoSj
bGEqY4f3I7nh89BmnYM8SdLRhUpJKg6erhaVF1bFhSPgpBwz30x5l0ellKUClm8s
HlSGMknaiOBcPg7zlADInJbDBCXUAxkg4P1ltjkO9GoSYp/ApgPTezj3tjsbP/Ip
pGzkjyssTB22u+NROvR4z/zmR+zGyNyn3ecTofDgsGb9b203hVFZfdOw6mEScr/n
JNB8rTQ3ofOHZTUW+fcVlVxV1UReTHYrrUxXwWKa59L3b+g7yzgRCCPVb+fcCSGp
NWTpBP1kYjp7noJLPbzO+IVy7C2yQYBbAIWctYmYnIOCbkDx64cgHJcbVnw3oaF8
IyH8mXn5QhwcJCOCNYMMcL5i4PQCLamtoJEpXyei/WIv+IJRKh9d4WEohTUAVOC+
dJeMvXy6luE7wx0VH7SZ6b68MURUiZVk0nT4deiEwQgSvLh/0p95bHOeRnZRXDaw
3EheCaMmFABt/mFjNCT8nWJRL0Lq7Fo+X0Et3KwEoe7rLq8dkY8oEs18xDoiMyII
dvkBe4RM4r9bXgkxiZ/kl430m3kunqAqR6psNZzkyZ2WNLxV4SD48oh6+yq1fVRm
yatgkP5eGIO86Sa0/XDpHdlyMEzKAx8H1cdRyz0WRI0jmfDTbVQEBBThmSWGzto5
+myrtboTsIvKCnvypHgl3D4kOhFVnDkw5fOQy+aO3wsJ91iUSQ6loqOf1Mwa/nOv
G6LMsUpQ25EYJK+8swUFEQNJJ6k2QDlCb1SHgMtpIZu3aQUKeQKi8lhkE6MN4C07
XeBFdza2axLeVcsgfhZSi97TANgcikGSSLzdsCZ7Ds0Nqac9aJTjcuLu8HDEvj7y
RUetkID47WXQJ0kadXWaZmBjHhD6YG/4+XIdth+Zjuenoj48gA9wF7VNsShIDiBE
YlTCLPb1prQLk58ceGoDDgfkcp6yftZjo3hfiJyehh3z3+E+EuQUuflpFj7+oitj
w8sbqNLaERGfb4ybTF/Q8V8Ru8UqnS8E/bwXVS7eakG7Qpc3HvsXgBvdzSNtRQPl
2muAPhPVCF7yCSzvZYBT5tBsK1JNI3eQKoPL9DpBp6z7iNoCwSQN/1NAqCvp5z4k
KqaKz01bqySbcvkBaX9ZiBq/vXpoWB0tZtSI36icVfxLZUP05kXO5CLuRmbQe4Ht
HgXmGYBHSBsyy9Gub/VMDw1KiDzS16fU6oLh3nZerYx+8wfBM24ThhluudiYi2KF
uupiZGTmllgQL/4wKIyRDZH0U+94qPIElMbhZuTPdfttgtL22H4HZjH2j1XDMxcn
XW9yZTrJ7+Qi1fC6GsUTxctqvTRL/b8lLuTKok1o4Dym2g0feyUUtjD7krU6+ZD3
mVQ8TGleXil3T8UbsdW1ciN8yUV8Ew9QDk9eMmcoIiT91k7Iw3kBU4KIuNXPWQpH
O8tXxFNFNrXYiMSpfFns1e9rcF4k8VpnDZvCfNpJSCORG0GGNVLq+pcVFadH9QTB
5HT8svTaNfjxThoMoyz0Zmqpd+ihyg8fArdqCMsU8qRkMDYjaQwaLh/H48cx0FYO
N/dieUfqPvfORQrdFNDA3MTvdbKYEeeDtFMOyaUlrQuopIMA4rP9ssHV8auZUbBO
hcI6A08dqwbAqjveI5x1Pd4xDdV6MWT7DEz89M4E2pHr8xZRJs1ll2U/CLl/ofoG
kUWil9yHKEGOF7thvQKMKUr3/7GvAkhNnSODJODBX2m+kqQfYw+c5HB8q9umg9fB
xXaNOHPLhY3MphSlYuTKJUKaA5hkYq9MTlWEARbaiGwtd/uXplN9GZHGei/32Kad
FN0olTcf/2ohLN3EXZZmyu4vk2HczQn4DaCchvOhbpwnFN0D66pd7O64lJtUbiou
Wg96skWAUEpJmuzFvJ4UwWZMr8S1ZZyLlOFxRiVWAGLU8xD8D/vqdY6wbgA4Rttu
aB5biNSyUfX3PaalVmZPooM5eOeojz1xoU00/4zG7aHswC5RbBsE2wghQkfUaoRW
5g9rqA+kRFBwrD3pWh2B6EgBQpGvnOanlwe6b709k5mi1JzXepiITYOs8yR4/Jao
kA10ttLSwj7Xe4WyPLOIcTo8/U07o8SzoK/72ynbEzHpjBfbu27NISGXx6Ck+Y/T
JUttWVdDPaI7l2+pIvj4Fv05lnFehu4oiYZYeEXo6VJ+M7eDEA4YnmvXRyNYx3wQ
GFojsScHZGI0dUZKOxe1KQvKhDgume2N0bbJnQmlWW3AoAI0+xRyiILs33GrVpl0
2gNvYrkOSGDon9M7FK2MYWLgtKVUV0dO9ZqNiDAzOfD+KuS4Sv1p8ed38CXotFrw
nbm8IMiThRePyWSYR+k4v9/niudBq6nTsOHdmnvGyEdnDtHtQmq4rVSV6ftCpbl8
fiO6TDY9m94ttyNgkkORq+tTT39i0mBqROAsyV2mNV0gl12XKAJIB+FkrYS8EGr5
QMJUVgNc/OCKLKQLbRar66InYmG9Y4RrNFKH20Dnu4v/eZgDpwsKZaieOjH/YWOy
AcMC0/ViVrrbJcjmRRt5X+LureLt3cz74uGXMEUmnaOAFmtq7llbwOJuLuT2XRm4
u3J1ETtJqbNA7u38E1AjzYiX9UIOxezAb4hyzzn9JT6bnkgRLjKtpZGYM+50PCFI
8K0ubb/WoerU6K3w2ynzmn6lp6JJBGqBDNirlY5zyfbX2jC+RmpvIDwMjBH4NL11
UUhbM0j96UKYajM+9XDWZm+qW9ONYX8nQkColFQWLvb7bTWJXdVDj7XFLZmbL3xP
FSY8ljRPTR5H8FnQI5gV6Ql4sS1n/0bnaYer/ZFB2QbXMxy5tpsLAevEqNgo/5/P
1pvuEMe0rkukPtEV91nwszbAhE7HSGqk4GCL4Bf+ChHlQ+LT7XdvuU/aqJg6Pt6E
4+kGTb9ZQ7MbKHzoxibmdRQ817oiug25xx8+k/gf/aryuI3Az1+q+EaibLIGqvT8
VKwj2LNvI7NFe9N78FwLPyA36fuwKW+fCUb27YUhBNkFPwJ27nk+jVQBMYrdu1fL
k7I0g9S+zUiQAZCf3LZiRduovnCQEdLEHGfUaaWCrJqkaMRCOC38nYvdHdnk6xtG
3I9x6WS7ayWAtlxbNCa6N65jlFnoogjnCmvdJDrkgNXdRuTbdO3ucWuEz7m22ZGD
G0Jub2rZHM/HtN0YRi/ietKGWP4pMYLlZA8VJqguUGPr6jIiHkYihUS5wRirv5TC
ih8cdXD7PiJqwoDxU7sTEpl3PtZOy8POTB743HEe4yLwnQj7ErfoBMA9usPfURGn
GNqM4IAz9AZsx1SQK4oonZNurwdSM7tg+wZM//CCcHx9QAmlwIbtTPXeZFlibTxo
5ugPq8+Mge9yriv8c8B6jNU4572HMlRXKQIAlOfjLWkO4UXw+l9+bpwTS7A8iFr/
akaeBG0vLWztk7TAuUSVpGubq1bcl692qrj+B4M8qCi2qE3LbUlf5M3rAAhoaP0h
FgHYEFeHQbmA9lz8YRUe+3Ebcj7U307fN+wq/OMrk8LodiszWM/ByvRemcaZd/3B
tRyX/l/eL6xzukCb590SvRdIu8ILIT6j1Lisflv8lL7rdFaubVmbt2mY1mYENrMp
/OOPEVfrcwZbhBd3hVpudlh4Bm2tnL1NId32gDOjJGukJDNYdpDFszpbTrftP9iX
zkkgzeM8ndjkyxRC/4RJW/E9PQSEnIXpdrBTuubvz/g+Nv3JavBiFQYFJfGefXDZ
xkV3Il3avZEkXP1kIfwtLQIORBNGBJ8aZsyzFnuq5SzB4gFOFc3QPwSu2Umo7XZQ
JK1jOpPlKEv+3lAvbGJZe/WD2wg8SKqQFpD7J+iacs8Sr15ZuPUoLSRUttCd3UD2
G92d+HDafO0GHrhj3unBxNBy8ObJVhZsmofMjnYc22qCEhEfOaKKfagyawmKBwDb
YlwyE4En53fDXVSXr6euS3yQ+g4GtnQrJAIe91N+C4+QnosysiGRc8c/V0JALbR8
XIjYzfJ/aIfVfkZ7jGPP4RaugIYmgC6xqrCLp72l39k0zXrUZ2o0kDI2fnyvWHTq
bE2JcWFgAajQSdImKvsg0EuvgOF1Y+XbtonLP9QkWhXCpAOVOCk73GqWnAsxonEc
8WBtEo6qWG6ohFwAQzIqx8kzYG6+8UeixDd5isPmr7iEk7mv/MuCFp5Vj9wUVgSt
/eSZos3lrZ2UfSOiPeNAJPUfCBKDXFc4f22uIKBEX5Qbbib+vhxRXH2SOW7FfPYC
7x4Bumrv+PNfMDdsS38Wu+RpqIXeY1e0VxQS54HE5ZgQNmM51B042ce7OYYamBA2
fsTRiwRqd3IMMtgx9My/xEi4rPPmropySe0ohMj4A3SMaZ4sT3dxNiTZSADa9izs
C3SLkijpqUq/bTKk635IRKkNJQjCbcyVogKjHRRu426UCjiwWBxVpbooC+6iEAIA
oK8sP4k81JaTQMyfS0K2yRsvS0IwQqKd3fGpLDKoUSlDTNhK/go4T67qYPsIB5fi
2goaLTcv3JYhg9+rHRUb4swFWLyyhVp/k2JThGWcm8n26FX+EMdki2VD4itWOswa
OJTNe4tEjHxJrYKPW8zXDS9ekyCV6EFBJYhXReXwxoMTyx+3KYu4A/RAm5OBqIiL
WjDpbTXvy00Kc95DqD84VSoh43FU03lfQDPhshy5Jr8L2g9V/RmvoQc0pU+gXEBF
wkGGgfGuvpH2kXrOUfcoWnT5RqBOyG8jyVdSOdv2L3AhGtJHklV1j35/bpmvrSzd
AcmzTFML9b2Jgp0GfVBfZlRmaKjA5EzroNjdNTt2JHYeCtVgXrpVBVJXcI3mpJ2l
QWgE/BcNyEaXeB1OfkVMi8FVC80RYLOcYNS3IlY0+kklNdxVrM3+MpwWErtsg+eB
dq5j7pcpT8Ly/gt39zWs7RqA1H7Prs2s5iCsKNzdTc2klo/9ORHYbVcrfDiXj6Ok
4mAlkZ84ThY2caHtd/8qH0zzq/J7TDHD4K2uaWa+VpkNxu3owakOY3q50q4BTu5V
vjqfQFvcZj6LGwP/gTo5fIFP9SG0U88SWlvjOvyWGdE5YN5w+yh+PpIywhXGUyWW
4zMf/gntlJe9h4wKg7GyI2jtfJIB1I7lZJbxIxeaL4koT+sYd7yiaV4pAPwoCBKk
GMpbIPAWE+lx+OJUlHts53DfhzLIDLqOC3pbQvXgAFC9DD3u8KJ5kektPgfCLOdD
iBy7j0a7gxmC7Hec1PyVareZ+7paqnPQ7GO05ict/WRrafh4Q+nIOmbkljxMx4VN
zfkIOz5+Z3Ofa1obOW0vHJUmW9V2HezaCdacLhVk07yVpwTBkLNls/XFDzc5zH/2
ZvIGf8KC0fDNknXZln1xdbo0hH6GZR5MZw4idxDbgdpnfK0fbVAW38brge2NGmrZ
rpBj0ti3VULfpN92nHPtiogux0/og4A/2gPfH+uwyR5VhOesKI9lDpBiA1ECWV6G
TNYM3mcOEuWistGs3YWQdJFSBAgWDpXiCRvDLsnzB1NPIBUFt0IdYWH8CtYDb3Ym
zlJCkFsjkR24erFIgGeqxPZQ0KUP+5dioabdbSm1OggrnQYMdpMfgXO+zCxOf8AP
+Th36+8Rt5xJuWzciiztv9Vo0m4amvXYq1IC3+2uS+3fcK8kozcOC9Gm4S2h5V4Z
aZRR6D9keKQNaVcicWQ2dalit6xq1M4cAJqG4X9cdHc5N246Q660zLFbEkx/wWDf
eNQJ5QLb4uLPvWlDy6ml0LeHfEyX/FFCFYac45LBGUw6YnVvQT6jA3lfeqcXc5pz
jIhTpU6U4uUjojIgAeAJdJztnTw8vSaj8VzjLMVj5cymQHb2ihrWk35V3prKpKh4
DoZjnvoybvL7JkbW8wbAsWYB/9eXjGkDkR7V4xNIQ1RqXyCRaiBClevIkQKS+6yy
G5uYDP7dKIAEzJ4vuNHVLg4lWNFswVJLh/MJGNIeQ4hYrKQLQiXfPtmN6IcBiEKO
Z7DpX9BueB/fSZmIMWw/8Hh145VIACat+WafwRayVfi8e8CAVFTLWb49xMjs6uz/
bVFyy8p9oqUN4XGqAeFDOCULyzI9XO4jrMlSZSXCDCwdhIhUjeAE/8UNo+O7kIku
gcg8bLFsvjVCcYm5EC9KnAHyAvON51O5XI+6OcsV2wejo4Pn6kUBmZQyBP+9bSWM
BLcMJdRU+iokC8EEIXzFpm3IV0peRfH5X3dU+9sdURXhV7dQgfzRLeYSWCLqjxHi
qezL1jHZQ9iTTTZcFNJW3Wx4AMs/RG7DwpTJX0W1ml1uThIApk1vgnquhFskR39j
4VSpHGhimwDTGgncC41os2q5bgyTOid9hiOzjl64HeOC2qkX1gcHgzCDVhKH993E
p0wAX+cxu8D2plO1VADioA6VkwHhQZDJI96DB34ItKghE+zpjXjMo5Bxm/LNf9IN
T0oYuhuTbvy7c9rtt55m04ob8JiIaIAAZ94tOxr6NMTGtCIgRGAoTzfnIQU26uuS
XhwBase2U5SFzCQbuN04iSnvdyI776BBOLXUvyK6rzWUyROr4fYe2mD5hFXJZAty
AjDeUiLICFYVncqB+eYUzGYLZLMZ0gxBws6YC3s1resD2HnwIVjJ6JRyTSaKHp3m
Uh0GS9TA7bFMB2eM5WdOEe8kcthQ/XxnGF5IWIwetXtB5vaZMShT5LC7geIgsfPU
K/qtieXwbVX0WtKSxdnxBo3ZfDswwdP9t8c5CQmqPN0F5I7EDEqgwTbrdyPLPaIw
PlsVo+NaGildYAVpHKpfd/Ghx9XjSzzdFzXdM+E0ji9sgHbNsKRsZUxg8JAgHMEq
H90hSUi11+87t+kJtQPoRcaZyOEODgOcHSZ49Lo34ro1S8Tv7wENco3unKR/nUuC
zH1lA+deI4EpkM6lwR3SEL7YArGqvrooRo+R5JHjEaSZaFqjAXl8v0z0RhssCPOY
6ZiACv471kJIKqknEYr/6REqW8bK2WtztfFiuWSun/dzEjcnYKAAPautAa4WAQ/z
TBfbxXdn921WZy45ppbcugOIcZsU5E3OWw/tkfg3iagqFIGwHnu5P0cgXuqkoAUI
JXjjDX+XhaqQO3GhGBTSK8ARYc8BUatApdt3cVIBEb1gZPDTApujFe871EwKw5hz
CiEkYCyWyFq8sC391E/IwdelHHm9QASt7323Bf9vyy0p79IRd9q8rh8soLmCnjWh
VjbqmCa6W/35DncJ90HVaId7dkN58/O5fnSiK26EoPqucwafCAk4COdcixJLMTq9
qiMxRmz6nKUjUx/FRvSy0wnwScgw7rpl+hDxuf8kjm/asnQpkua+WhVJDqDtx+PR
ftj1ZhCzgrzFzc2Ef6lnNqJQrfmT5Lb1K8u6yMCI00CEgbcAC+sEVli/HzngdJTW
TdlRzBxQwdL018CoYBfddGdjYcvGZcrtx043BhaLRR04GCWqVn65VM8aw+PhcsrO
OVPYdSS4J5vC4vr3e35zlGL/xryeUiBb7Dt8AltiZ7GBdCK+2499UpRNmOBI8Q1q
wb76ANpmbnwD9NPL/Me6Hzm91yFKVG7O0PoCGgTvw2RnvHrwLY4yMGYlHP3mDrIK
laSbKKSGGlybekA2oMCe9iiicStQ9Ug9LuqSeEUX2iUucWrY+TNpWc5nlSwObbIm
wTeynieqKmZY5In77wibWCSze/SVB6nLDldCEDwrUfiZTxKO6TOHGYR5P6DtXyER
sMEXMD04NqC+Mgg+LCaw1/BPThuP26pbO7BPya/O9mWSSjanLx8Tx8Du06zBckyK
mab45/1p6zKt1yF0P7b960MGseck/rDaI4XNUUs7Wcs=
`pragma protect end_protected
