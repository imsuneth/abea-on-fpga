// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:50 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
It7a4hGFMqCRcX9kFcypujEi49V0mALMS/VrvnjLA5ctLBw92gmV/52bzLA/HJAV
HkHKmtDFudxx5sN3cgxOLtMytmFhUNEbWyA4jXFJIz5v0Ny0o0Vj/D/ThFfNMoPn
h0gHnk51V7TfFGLCI8j2X00HaUXUoskZJlYEu4YC7XU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16624)
piQmH34fsZLGqeZib8v0aW5rJPjWeAx6NySFm/cGB5Qto4jc26t3G0fDuW0zcAm3
CPy8n9dTsb4+jmUji9VEffW9KLhvy0dJVwlJp2rOSNLxK6mm/hFEK7iWxdTonDgm
4NXdjekQIVI3YGNo8sZeon3QOofzX3Y42EhEl7QXsea4/rzSfpezag3MGaQ3Wr21
PrW7giEDJGOWwLoPofzvrGUTaS+C6lyI3gwH0dVB5C9T2TkAO5GlZWMky3iHMyXn
OyzgOmhN4bpX+33Icyqv93MQuKRdDoIbuStrs6iDGmoCACMBRK9t+wVVM1sGiOc3
Uad6Ci/QHRyJfSTZSdpGH14XknAsWlXGmOp7H4mHlba2+fQoklo/r2DtIh5ztUyb
B1lf7bz/BNK5UFNNdzFg+Q255OaYoKIUeBKnu9R7pirCZmixQRllUOEdZY0k7LtZ
QMrQNwGkbGsRYcSZQAWMmpZP8EJwhU4ifoLG5VpuFZMUqd4mJNTd4Ai2CasPQtYu
sptHIBvcBYwGQkgwc/pE6t3HlvtoxbEqBIBIbdnHnWuuqCOXGlkr5j0aGX1eLlbH
iCM8Kx0ns+aALtBqvNea2V8V5b/wimGOJPSWPpo9vNSkLR/bHnEIf5qltkI0XCYC
zL0Mag6iTyATrReslack0MEWiJjDXZCGlC+VxUK/aNln/aJza83mvcbeFKhAW25E
rM5FeNlymrukzQGCQhIrfhoqwxWryb+SQehCBm79sztcr5hX8/KOK1Qr0jG4MMBF
Tu04krGgpaznTPyeK9gjeHHF/MeXLQBdLiG79zV9aQLjvud4ZsuHCujtKnii4E2+
IXZPAhueFhhPgGyQEuqKzzjaLM+Q/P477pavfCKFbzCU94FFnmw1gXGrGUmShSI2
i2uY1htaZckBCL0stJXujuLIXxHEgPv6epCjBPAqpLmDv7Zu12lprPEqRqacqic3
AX8tRl5gUf6GyByBsqd9vK4t8MDEUwW2JgXK0xjMQTZ1USR2vVBoZ6PUWGsmVHjn
mmoeENZTZ4a1Kv9RG/vq3Uy26tzTtYHl4WCSAvr2hOSK1cKW/lxTBdE8ZNaKwQ8l
B/6uq568tFHoyPl3wxdONY7Deuc/WgRXgD5Lc6q4iKROphKKNwuK75LZaPEZtf4V
QXAij2aRs3aHuWb/z3+LPJ8EuaabUTUyMUtTEWpGu/HUmZmM17NGx2M5N8mRMS/z
pQq0gzMar5e++EAMznO7iMfHLiZAA27qLOeGjuXVDWv0cuZEcDQOHsqWDpdA1He2
pHTaBFB4x4zppruYKFDfzdujIObepF94p7m89FFzyl8AYSsbL0v4IzDLa6x5zWo2
43ypH0dP/LG0ATY5nqKdamdWTDOsSx6Whef96gS4crrhzK8edKHmd8Bmy0EcNtr6
M9pbN0be0BOr0/3Kv/wIp5g+gF/NVt/4rQlVXfCYmqDNFirvTDl00S5TtIirlTnU
2Ezk0YkkscBX2Go3KW2LLSZpt+eM3L5kxFrkdsNMiSNFro1530fhyblE99Yv0ZAC
BNmsYJPmqebsz4nkt3sZfec+VWMEvyfgvPMKAlkF0jSBfrl62/Co3fcgU6I4MLu+
UI66rC8kZpLhdO4jFXrXZ4+C7BDaVDZrx5QUgmgi3vtPEtOGVboydmB7of1SFdyQ
5sCe34HF8XgSB8362mPP0OnTnKdKgUmWdw6HKkZRrIPDopBaI/kvF7awTSH7WOzo
JlpAtgVZhmf3nODlL66Z3l89Ze2JJkQZm/WkT3qFZuOpCODoduAlqkyFcezPJdIb
qkvDASrbvCyuO+Rzvch6V9yPAmMpuX7a2WQis90XPpfU/zylcrKwXYSSSitlqBIV
r1flZAuc9TNp/Vx7A0+sxqRJGZg8tgfMRGWOifAPVQtnUKKezf3COQLkuLhT3wlX
ZhELl1aW9TWt5sKtNEKcd+RkZqn/aWyX2MCE1pPEdmHGrmvzaSasiR7V6a9g+JZI
Cw+i2118Mu+mUdxKsd8D7V+cMbXQxuOXO4VjKXqbHTitXH04ZOtzZs3soXrMzUz6
Ii8kwTS6Umd5Y3xUhjqUwjlZfE7VyKpt8xCbzBIR3R2hYSPb4fd4EG9DMs2Gq3hi
KRxG3HmtHWDNXmGH6kLFxRVp9HZr5CFCVnLqJ9FzpLwMaAFvRbFqbZ0vTCwI1B4x
Yeo4wkBSrKDz2IUIX1mihUAoeTh82UKzbWrsn0m7xb5VG10UciNSrtCULhpqWvHP
UFXf1KkjG4DUc6RKGmeN5k+A9vFeeG8H7EgptmMD6e6Xqw3tjaZOPDPZaHGlrJCg
lTVNrKUXxNOipHKbbgRzm1RxLInGVrRFdUxOskE0cLVWMBFxU8OdTrgyaDf1mNjl
Pp1mrWql2xfeOXjwfVbrWCaaGYNFxvSb2uIlLbA4vtrU6SicTdBjdS8AxxwQu8jn
G0ITKa4PDxy0MNG9Sf0XdWxD/aF8ww35iDjG9D9jBPVBUZiVxYXnMOyIC9aXC+V4
2duW5OJ5hpcRrnx+oGCmdiM0bt5ogLokqBjxo85SaRnyQcPN5xYkjBsW9ozyVHit
ReY/0x9/GhtpDjfvptoP58GwBTrN0cvGTEVOLxPFux8fHcjIIMn1Us3/sozDUwWr
ZCR2HWKz8RnAngN3l4H02A+mVbGQhpbog2M9sC3Ub6hvhpKhJ5iemmP057ErRU3F
SdpohgP2F6e4SOM4L44TpOtrnRk+xySQAmO0HHwTSqWxr7ztpfIDljx+WMcXd82v
OES4fg7ZQYF+KPzvZW9sbshYns4VsDB+L2Lcr595CFzR2J0C6mY7mCxV4ewHIf0J
+x0O30RNlwcZqvT8qtzKvVECyWaDPFEKFtbFYwi8NCUKS88HPPaYRbrIzRQjfTSN
2opY18jmLbvAY9cZC1nt4SRodIGU0n7kXY0Aleq6acdY/aEXBt55bb1Jh0s9Y9Qs
G6GG2NuS0e+csD67+cgLuH4+h+PJJhPxl2Il1Tm/q4BgSjr51+VuiFrXnD/+MjZq
ciBnmCgmVy2MPP+NXyXLX+xiBRX4sWYO2aqpTi7kHXl2z49FUvOfLCiGxaByHsUO
GhlQ1ClNZ/1/plzCLzOZ7+uxpXrKBNtmyTFuL/Q2j3VwWsaCwsntkjc9W9uv/S10
JFk4pvBfaL0i4D4GHNBNSKpKU4Qw5BMLL3Qsp1D+pG/vAtsQO1pmCL4vyb2PW9Uu
6+FUyc13s4mfew/0kgpj+LPZXyXVh1dosQYyeTfLGmczrFPuyENy1Kp0kLFnoB+A
53ycXRDuGJuiLG4A914sJQnuaxmqSURq2eRTczrc6NU1XeTe3yrMzlUtmVMXzeyi
WwY6ZGtzThPA5LwxVASxCdoHdrmTZ81FsYVb34regzscniTvu31lPbvWIIkMBSbW
NTKLggFUSxvwNwD4onQ0sMTIPqYaIUgKPF1Khw0YeNf9C4Q4dpZqCZ22FHKZmqXo
XNAPJAAVZUJ0WkVORuoE9EyqpW4G7QcfxXc1t6RbBo6FTPCxdHPk0O2I+5XfF3vx
h9n/XL1NrjARJDFP4PlaUd6qLCTNnU6eqLXw23oqfW8knLgi8tPtSpbblWDDrTgs
KBjzBapOwsfvNX5PSwQ98i9J8IO/QFbQxLQgbmzvhJWlhVGWnVhHZJbjSPB/MuyS
Zo4fF4y/XErotaJmEyhpT7y2X4wa+LYFsTCv/Sx0qoUXptZFX3o/HRKCTajucNan
R6Utl1AIOhs4FSEkuAGarRnTaz6pnASELK0ED3ccy7ftolBTi9M0wucH80i1IJYv
U6HTCTadDOg2o4JrdxWa/OeiJ1DFjyOGpO1GuOV/Yaj+7gKZlumHp4pWb67tKeM5
vCll2LX1mdba+kSmlChYYklrzf/nElL0RMsix+h9vdvIPkVdn0/4nz0lubL+X4ac
KpShar4UY7/LYdbc+dBk2aPfTsqzfgGE3zPZSZD5Ot+B3ENTihmHwbzWC8p2J+/G
YR+9DUFmWhq84TQQSuTCvXuapqtjWMXioEUWvPirCsx8a4sc7N8Tu3y9HAph5ZR7
uRbIeAafAdaVI8DCOw7pUn39uaYqbb0MESmXoK8SD6+/rj8G8Q+ndNB2Zfmg8aUP
gm/UxGI1Bb0jHUz7WagpuIQBHHgaru5XDRRPQSzNP7M0BJQATgy4YoaUSLcojVvL
SK9LJS60RRJ5hDP529W3Ni8a9ytn13RW1ndtQufLtbga/lAAz/jOKZw0PjwFgZsb
57+T2ZA1NGzbyzdt06osz8zw2/gctxK3Z0B28VmCZDcGzTIlmWKfDFkdGRKBvye5
GheuZf1UFQpymcg5KQTQ9K/aDhonVJ4ymFcuEljfjAPyKMn5hGCJ44CujQk1cWHe
LDnwd/X1ftPCMCX0QqMgIDM7EJWK3P3NASrjl1DZbk0bFae0sgkeXaMwnYRJ5NBb
DhTkYAvlLMZv4nvjNpjMDdAAKvF1o6Mq1p3LApprqRq7TL+J6LjYX2Ss/CtwUwyr
V66hs/u344oHbL+OtRfdrH3TVkZg3XJPD9+IAFhrHsrB0si2soT9WuFPayzZn6EM
vx1t+WPnhcNIjRtXz9ahsejFgip8BZ9mbG82wsEA3f61ENQDlszPql2tQZMrBF7U
5eifNdVTJBtLq8yIZEZStwHUtq7dwgDj4hId/X6J+zXuEexZdFaroUsiGcQlJTod
1hzrLULfDvwAex3+mfKyRIXjyz6JJlJY2r830JEeTwNyZp6jHn2GWICsY+4Rfno4
y4UAXe6WP7vnjOa+9DIrfkocenhh8UQUlMTiDh+8vq2QZi4UX5i36LORmgojTVau
eiKYW0ey+rQCkf2PG7B7oLN4wh1R8oumXYl+Mj2RQ0IixfsrT8wlMgH6npHby25C
2Nilk3+cZtS2ZxQFANV1ypdoU+9fuvUyp0gAP7uuj9eEG9AFzIfUE4Ie/66gzNTx
Z/YMVIVWSDSIgyAMvH7CXhVL6iORdyZGoYB4K1WsOIiEyTxrNVyILCQl+59zP1si
OwGBFjUmPf1I6BTEFRQho5pf0Zs0RHeJwQ4A5iQxmiZKXuoqaeCwgPlSCTWVV/oX
Rswn8IFrjo5qRgRHU25KF2OvzIpRM0ChY4DTSxQ+Zsjvqh6J6eKdvkcv5FB2Rozd
pUWtomn6CTNUmoCaiGtypJYPQ6PmJaoH/6eyrknoRsn/qr/xo8vndKok25lWZG5c
RKWj/CytHcHBd0Z+lsbJm2ymI2Ga2ktE09cuortmvbqs5pEek4140xUlSL9e31PB
yjD2/gEIvClsjNPqCfhX/S2JyfficpS2JLVDKTG4SXde1bISd1oQ3nsgueK2gluh
f2qoSc0McYqBquav3A23Ir8INZRoRV7bz1AfTV3nZ2cDbODfRHDjXkeRo2URc1rt
CYafsmDSDJC9PxklIurvqk4WujqBXj9ZSQ3vIdCyOBx+94HB0cU1nZaZvyoIacnp
Rl6qTIb6goms95LQtkv3RxyAsh/MBaDmZ7dYxPFbZ+/1qZZuuyJJOou1XFGvQLji
hUh2hmyWLgA/LaphDTTBVsVwfXsOeub05X0QUkFKJ1tMEBwMS/+Z35MrYla2rDFk
1AjihnZADyZVrKAcAIzMfE6FBBW5HIIiHsgikzpoWFPSCB0ODmKGaLtked+o4Azy
WQiFGkpWgeUtFw+HSYtyTRi2VTH1GsBG4Jz/LEXBADE55xCvksmQ031D8zMyVE5t
0GhA81HP7sAmlqD0m1VeNkZtWWg6ibecdDm1+SIm+9hPEhznMAX84pUKKlnr8qvd
CQuSfIN3pNdhN1UYpC3wxXT6VGAOLmiGmBsbmiEBEheciK1CNxssgcglV9CkhWIL
llfhAHdHF8Sv1tF4n+t20LdU+GWFkZ1HtezJphPJLtKhtpS25jSojkJVHgk5sFEo
1ZuKyYwfZCxbzzg9ViETbR1cF7lsRleXMaBR4lBWy1sy/zM1jGbBkAyVrVaJSUKa
cw8MILVVCDG6okVGsDIbAJfnv5JeWiMAootMmf1nM736q8Wlm/mjYvEV7eKxu1T8
CbpQOlWaP3d0j7CNi6oyLW079RaqayutFmVI4gt2PYtBFfcUuqmFgIIIxUOJ/s9v
IuBWPtt/Zh1xYdEQsyrDfa1RSUE7+pM263IzK+++jKP+agYr8TEBVfqTG1n0Bf1b
KZvIjtxnF6XlEsxakVyPdrEHXC9Xi1IjW/kut20hmi2kOqEExoIsiKTotcXWYNOS
1ujshPtha1n4yYhUIT27duMRB6kfKb3AiWeSARhMZM14mTrC+31ut2N0F/njEwst
rQJEPsOYZ9c9GBmFt1E+RTVPDWKgQzWwk1HKQPZle6voFfq0d1H+788ntShNkuYZ
MxnEKcaIiFL4RLrqWfS2R/CthBwsz44a6LcLbj8V+/CYWbfycJ+eWXX3I5DyXPJg
/lWZswBZXhHzfKg+dedSymYbnXLIZvYTPy46Oo4IuBkOy0te5pjgMhyV20xwTo80
DF63Zk86UZUoTici58yUmMVv3cz42CMJBRILxop5XtpJJnPK5GeyNIjjPjf/FSJ5
1whlRQ/l+VIqEnvAWnUODQUFmbZJMyphQFzErxhsUAD843qP/5X1v51ZB6X0Uet3
WIDU2Ryzc2ebFfzxqsWGz6J+2p+woa/qwPUmI8LjYgymx3ErY78IHIm+1xO7IXS6
E6t+iz2aAlhXme4tDkyd/La+pKGD90GdifkStTYujqvhTU0qvE80Jby67ixOCgeZ
4WYhmbeAc3nStdnCNkXPXNMnEfqG9qkbkPoffBoq63cDjocWXYwpB9Kxv0fqQeKl
xpj9nG1v9TvqCglCG6IBouXdKS0XTJKupGZSqIRgOuvuy0T9zKL/+BZe3BVvLjQ8
ry9gaOY/RkEdnyHscp5W9wOax1EJd1zFjKstpC15CGnllbJSw0L6CpEhpgIk3WoG
Jazs1G74FcFKZegdEUdZH1cvIvOaYr337lMgvebHakPmPuJjq4QA+FQr/hhUVysJ
01tBNMsNqZDHiGLgXsuCOObLsckTZAZB5pf2asQhBOpDB0D4C6trpviIBuHaqrLH
VD3AKWNS7kd6KtTvRnZFsksKD+munAZ1y3DKfXe4hKMpNHZGo3Q8p5sE9vGPW+Fh
Vs815DI3DvnVC84lhI2r7ijd4ubH1th8k1tNmWCFMlT6jnKmbJT3i43W01SXVIo5
TYO7attzsKUfUiJ8PSklDXpxHUB9cli++WL+viwll4fuXyIYb9903e9sRUtG0jOX
JYMOHhJsiAMBRfUORi1KX+mlCyJzHUjorlDzq69pMXbJWffik8ZoluOoFTQXlVit
i4V/gVA/y2s9V1BqxKJ8WPHb3oYgKVjg5GQlnNDAbEKH9lvEtue/Fdp7UWQQ1VfR
cGwc1k0TuAXchfZ3aedAmbziQbCk+fwOqhsIbphBUoe3ibDdXJXVtlo8Vgb9ImL5
b+C1qvfHB37ZTPJWkZU5ZmSDL2nK5aVMLYdOqulc5VVCfiMDQtKTK1WOMq7kynCw
V9oQdxIprtcFtKMXVgbjUx2FxpVzZfAXrobNtIr3NUWaCQSta5FjNMDkqxTeax2N
xe9ZkGxgrCkYcB5QymIiqTTFY/yTOsunzPY7iZaayzxpr67KSHqZwDYz3H/c4esM
hLSiFM3Z/mdQ7MpASOh6o9dlwYIH4cZtVAJk4lSypOrGa7orx2zwi/s3lM2DHBH/
UXK/ux7lZgsDEC2kzK5ASWFuyWAcFfY0GwGqGNfs8IP6V7RbVg6mossRVtz+YHO5
hKBMD16MddVhyjwX2YlJkXnQhYxqEJ1tRGxB/N7Y5CqM9jrzU36Ub8iBX+pruifv
mTzRYSfxlh1MNcr8o9MKtf+5XauwRSt1QpVbOet1rhEvy4AubfY5CjCfuT3NR1c5
ZFZEuPFDmvCySs1TE8ZSFDxyHz0ntspVeSioIUOgUFOZSxCJV+ofmPigq/X0qUT+
cOaRm3VpX9861svynkjgi53ZcBSw54+JW+e8BtloCiX46Iw8Dt0qvzWd4MZ1aXY+
Eh8/y/jMjYQbJvxtmjgkqI5eAH+uDmT0yEremBXKmWIYQ2MPumVtYLkglD0kQKO4
yYq85SEr/G7lOdKUoACCeMr+tpUynSCBvKfgb833jPmWs+BpMiE+wDAM0nZC5rhT
+wo7xys4PRnRAPAlTT6KRtVf1oeZdccqCp/2q4WRnQZU1Of1ay/XbnciFZqCRnNd
Ya7GZR7g5jowyCnLbKUpSTsmJsPn+1jRSaYz5slBKEwyn/kU1u1GRfX6IHLQENLR
+thM74b+LUSpIFyDctYG/2BLwSvWRmyww23UvVNfHrBlf0/K2kM2K1M0ShwN8qQC
CcvfKETpSljCasx77LiDSVafQ3OA9eP4epcX4WwwLfFZi9X4NXWaw/d2C5ZY8Kfy
LxJPkqa9qmCR/CHGCJshzmKWRfac4NiUo6CIE+tXkTGN+gYRzvjBjPCRs/pYxsoa
nbaupM0/sPwv3wvRqIA6rjX68che9azvX9kF1bxAnOu4lSQ0AcI92nirYOXDbLdZ
t5rhnf+epftYnF3MQ/tOeV+AAy4bWxQWP5APF73UiYW9k3teB6eTjMn5lBOvPQit
snJTkqbIIuc4dvzbDCsd49gftY1sp5fqk4Ccp4nc6kiAut1rcouBrlSDV31zASKP
hx9TWc7Q1AQJokJQ1WvOuzO52NxPH7gd6GLSPworfJUK+kKw8WGiI8+Wd1CroYJl
CejJwIqb6E+oShQuRFBo8V3I3j6ul6vTzktpiRJoTJV911KErNSK3vck+LkkRpNd
oSVac9OkfzPLIEAo8Fjtm+Z8am7m8hL08/H2J0IhhUFf+F0OKUKug6rovsamNQtq
8SHzYxtAmYBsFlYL3GOJ5m4aeBnD59xaaM21FXUZMEbCD9PAnMbEP0RAHxCa4fv0
4dbLn5KilsC3C/TXodQFuJXp5vXKugcooPQ+LhoNtl8whRsgMxzRvT8KOT8YXZUD
ylugKiUWJ/+kk3y3Dj9HoLY0AhgxRzi3Ef7BLxDRY3PmQQ+6+c0htlhYS5aPmwSX
gGlaxQGw0VW8DTePbo8AD85e7tthh3bBWSvkum2WJWkgnU2H1lVKMWiLASPDndeL
Qf6tJPWOBnkBwnJzmA9G0t48P261+86DrvC1lyj0GLDR04GnXxefMqmGoREF9OWf
F5qlPN68lxYSxauAk32uEFoLUoMVZkHpB1e8a4EFRj7Isod3/+VbtBZZcHzr0TTP
eH+ISBV4HYpAAw3UVfMxv1D5OL0Yn5K0tfhiCKB3nX0tIffuZNcC/+CVPbFLyDv6
/nbCc49/fVJ4koB4AYk04Jh8/BMl8fiSLQd1tn6S4ocnemcol0vYTXDgW4aWu/pB
MsXBJdjVmj6LSvGpueEG63xc0FPmS0DYUm/jKiKzUry959lcg8nq+KLms7nKjp5T
alRYKGI0UN6q5VtlM0rizaQ4nGLLm0G1oaDIJrbo4Irv7XlGeMdY4T8z6MuhlVtz
5CBLsFPHIPyK8cGmPKtAR4vbSsN0oIUbT3vF6Nm0HZC48UqT4IT1gyFRE+Ys0AqS
IJlusT16pXbP+WcBVJVJ9mdrkekncuTzvC+QaFY+VsC9bTB8dScobCMl7VFp1wLn
cB2NvenOqqoyAHwZ5v+ZOWChD0BvLZ0GYbQASWvRgQZW7ISSn8YxGuMjSLudaesY
ZMeEQ0c2G1sBByv/sbrMneXYpOv/vF/A8sbJ5ZH5GY88ZNQkk+9cK35Vrw3hYmNA
3LTeOD9nK0IG2ZPQFnQ0CW1PmzgiU4SabUwCqYZEUrpf8qV5ZJZ5Bn2U6svz4FSh
IQ8TJVUU45bb0bnwWqT+nvX7qa9hZ3/TQCCey/xXVfhmBrPvjHGri9U4uXIcgIOq
GQUbOpru/cvM/I3yDr12eQMgarArewQG3DRsL8+d7h2s0yaH/pJXMuLoLIqx0/xD
xRkCtci6bJLRMdi9OujVS9r1o7NIEq1wS37yybP5Zv4HMJgYMZLP89Mal5Cht1I8
tcMsuC0beOGpqoekMN+fDRFtx/5lo0J25LTNsPp0EFXg7TXYOu57S7FouzMgtlao
9h/xnBaQGDKuc1pVTrRydbcIcClcbIkIUcMVBTI6YXdkJfhWmkE285mdUATw57EB
G5UiMYoezDQukEVCJEaWPLi0EmSMPAFL+Kk9M7qxoQW1CCPtQnpHkBlas3OjR5ns
ZTkn8IqX8HGMHFaNrvBBiILSm+szhqVGqPkRDTFkJLYcBFM7gtlz8jGMw+FXFB9c
WVdysCKDPsPBIIFXUKCgo6IYFEfa5OqcPW+A2XtiEGbgGWk9u+4T5p39j7SHW/Yc
Ab16dUwvAYAp1vSvb4/9nN/bAdhRWIJQDg44PsxU5eOpl9p3ZBRvKjLHnTBpQkWq
d9wAFxxNvy2CWtBp6qqsRz/IE1GQvxJq2bYWzL6qTJZsB1uy+fQVo5ObShVoS67Q
K53nP9LYIlU8x81dJ/7Qt/ZUgFqCQCD3ksiigbSaGKRFQvYt5Ry3uwTfDPd0/OJ9
iroI61TE7Hj3g6BisJ0eShlL/QB4RT02E2eyFH2zo6eAIdvaTmJYaZrlvGyqJ5Wl
9MloUeYt7+8Bc5Wd5RuLnAs/kTZ+SW9+d/NMAOT6dU2XUzRfvIZEuQ/whu3ha38E
spkdpDTw/qAmxrpCTAScsf18JQLPFwsw32LemxceI7VUETq9NiFuW05VBUbpoBlA
jHsAPhWV4Xgkw1Kt58hpIhrYx29hfjNozJ5/8/gHQubfS+TeZH8jw41vhc1vln//
fEXfLhJeiQnFPCMhVB2p0b1n+RloUG0MEcYpYYV/3IcwTjy7osKHZzJXvaPICICu
LRP94zM4tqmCPJqosolRyBc6Lpd5nVae93OF/kLtHwzwuMoowgE7+R9aHpMfv9Iw
WsSfl6ScO3ulyuSPMk65WCaZ9JBxLzdgcf8hEhkbenLDkX93AOd4/Xvq6b4/QrWr
qzlyFnICLVTXUlw61R9tNETCiy6j8oBIRhcei9q6WxP0zt5Hmb0wQWGdbJoqNsH5
yhPu9r4SR0S7y/7QGkGF6623W/sgbheifR5GytGG4uuHVw3RXD+2P3VZs82nOqQF
ha9qjB26T8wDYnjlYIYkc27c0ZmPPot6w/IIuWF+BwGM7k4+0svYwQFSqNK+MTG0
mrx+ifJLHx+1cTLScmMSOTRHyRQEb1f+I4tkibfo6fZVlTSjae6V6X5I81TprKKk
tXpWpLlOh4KCk15iWM7z4vyqVxbz+K48w9SkaX8hXFflEFEQ4sZYNtNxx+vD7J61
AYeFmZkX1yZt4Oj19zU+f1C4cwhmMZGOhZUlv8devgIT/XySGb8w1oWW4G3i5Hst
MOEcLcP3Gvjx2VbEIda6b70aaxdANoABCh+8S4xOWH7HseO2G1m6tKHF/Mu3PjgC
TxV3yDH3CgGT8PDDnGwzyhVJRXAkRBVL9cSW6xmqfqM/jJtGtOAE9DtNAhhkIH4g
Ou7YhMoK67ClLQVl/K9W2BhXRQCjcsJLY+7q8yHCQwkW+MBxBCx+/y0LbunTzstC
ZZoIhJRmzES32V40Syi67GLEdIetMjXCkq9LrtCpK/+A397opEcFcxm61yvV5daG
bW4IGGSG8VM0mLAQyPbdN6d8RneDHxC/5MsOtjlE21DktXNqaq2Fqua+fYlPwyRA
CIkOWvpYG/scfcCAvXgguPLDEiMU5ARjJrYQNg2FRZGnBGNaJOXQpohvYvN85DIE
oEX6/sA+u7FJJfjHuYkPDI/MLb/uTyOFviFc2EgpITMyqaDNFaEr30wrWGHTf7zV
QHbLcwbxbEyT1+/as9kueE8L28gewkdWOUmWOsU950PAlyblX+JYvjHphQ22h50E
1+vjvkwx0FZRoqVFcjBtiN/X8HBXdjOJvgUDDaTCsst7QGLBaP+xXs225FX4gh7z
tR6x8gD+PkMNN5K26U/qcfqVSiseQLyRpokFVhEVSIZ4VPGK5o4K8gmgJ4BN/1Gc
K+dcMqSqjvEJdPOCgLPpGLXuWm5jgyIDmW8RSMq8MyOJnKNAys64kaSRBvKe8GwZ
4W6ET0GktuUhqC5R4zgBbeNbAYtUGUs1NFkBY8vuaM05zkRqSqkzYEz6UwMcm7Ig
w6XQ731H++0E2H4PKLS5YTpKU+xEphoToiKnHvbqSF5XB0h3gVBkOoyXU75zG+HW
+0xj5LnWzGa2EuIJeXv6eGqiRXNe1KS+bKBSOozwjwNtXPwIHTnSRKF+fng0BgmS
IBVqeZ/ZtenB310+MXeorw/bRewfNiz1ng2yDaF6sMbNR3LVATpxc2/rPGkLhnXn
Pv4bUobhJmB3WL88Mo1zj4QBEd7XkTYgDTFda3e6o60VPqhlayqKaxiXBL4KfErU
ey54g+8n+pfWcXIAAqhJBlGgISD13/ON5JERuBELZdI74kBBjNOqLc0TQQDabkcg
jGVKNrUqLCd96ZnRkw3kXLKvnoHcs/SB1YqXtJ/6sNzn821WZmAnfVAo+L1z4IVa
micKh0hywkFupGiciuEqVnhc7lnjToUWJJHgOP4p7iOwQQfhYQdFICd3LwQZuD4v
kKLN/GWcfcaa5czv4PzUM4tnkAv4HN33fYJgNb0c7zOn7P2AtsUQN+vwhmn6jiEI
oJQuhMzQ3zWhvD53U4BxTBriruos2xSesM5ZXpTlVrs1/Z8sq41ZqDOFUSgR0DdP
VUkDU7CCJSb5ga9bKPtFBnO0BcIdoLVDHP2GmPQXoWZ7YbzVRW2mrYxyYpooekks
0WjUhWy8ojarcLUqQ9txnV8Qk40R/pssw7kxvPIhGrcGajgV8ztfWRIJ3Um8RB6b
/oE6qQ7TfLdpD2VXG2kOlcO5x0OeWzF5Mq/QxPk+UryvuM0MbDdW2P/ba0YttluN
aq7b12sovD+xpADAIrCBu2rmf29mESDSgw7aeaPUb0cX7MqGUhFhirzpRyLj/EBj
TYR+ngy97KXYKjrZIfVosPRr5hsi3Z1MkB5zo7BjS3Z29SdEbFp8nDDMuMd054As
UoEzkHvjEfoKfB5cJ5dZzmfGH0MFzZirih/lNKcIPqAPSkqHmY3Gca1xwN12Whkm
HNcTGVRUmiPNseqTWhCTBvbqh7D1GMmkv3Dv9PmsBAxeKf3qHskbB8BJKp0gcx8u
dETCGTqIqxxE6Qwlvm7H2HuuOGK3h77wDtZXiMi2YlILSDFqo2w6TwWS+JXltvF4
nW9oZAq0arDM/kpTzUXIWTlNK+/CpryN30/wAt7jx0W8Obu1juLz3EsIY9/Ze6UM
MlRCxtvbMKwVPIWSlU8lYIPvMzLQBbUsa3le8nkqB6pVYSeASTXXFu6qbmI+A2Ql
rlVDQzgYUBsI6pb745vDZI7g0WNZVecoZkxzAh+twAeXyghbZeZ1qAgFA7ng5vWk
pOhFk/if4ocoJixS7PAJsFxffkDRI7C9tsa9vWOImPicZxVZHLzFtT9J/fsqy0Im
Zhd2sKC5F8NKvJ2BOq2SujbxGVmSi+/y85bZFt07Z5kt4p19BDmyby0z/YMoMmfA
rDyfxC+hzhKFRWAXRhdWpBfWP8j8gsp9tFm4Mcv854+GDp8xEwuA7tivtW0aWS/I
d/wGOxkl0XTCF88Em7Fd7N0W6Nz7BYRPoYFW9+/jhnzS3bId/QZiWcodHNkX/UR9
aIwQf+zSjR1UgV58r12F53rBx4h7/2InCJM+E5uHxjj7C6n+kDZ+5qeQa9dIWRZn
DxsC6UJMLx660/LnFQrLwEWIYFxDzjqnKnySEvWja+7KunMfcpAfMBNO4xPL+Xst
uJlgOOTMlAl3uzETKaO1GzKDX+tQ7hBkMuciiVuQ+66hQMV30oMrWk5uB3eC7vAi
wRFezBMyCI4dEO6HWuFMtrplryo7c8xV8wWU/KhJEZFOU24HPYgtSztFN4n8L9kB
f7g5FdkvRH0YTQyP1r4c5Fu2PVhOazYZcYWNw4WaTrf83zd82Cx+FJ/FuOeaDXov
3zGnGY6cHXydV0qOghbm4azMqiNj/tOY5ZKohH4qUz//O73uXLtm7ANvH0fsZ13M
FwC/KBWrifnVIpjIFK95dB13UplmxNUnpiU21cMYyCzChIH5taibMeEoSYkkBZ68
/j7RcyTafAifiP5ocYZ2YemHQWpu1DaXWLKrrwZOl0dU+3PS4qKn6U62oe45ogm/
2isV+G+kurxBqtAAZiNZ0azr3HH9ZhyJTAG1wbVfjnfag4tb/yvEEJCF5FgIcPsS
vKFq4FBoWS8AH1G2LHK6uf1zbX7IOtiX+u9VO2FB/CPJSy7821ZOsnbq9jrIgqM1
Z8TjKOQV52nfya+CxRgDr5V6Hc9tQO60TmwZKST7WgxzbPYOcJm9/lQmUkJbOXRR
35NtpELNkRjcL8r+kyl1WzwRXUNzYhT5Ruv65a5ksvvBdZQI7Qw5rfojT/spIL1D
FMTs0tSukLQ1ORVfE94q61ZuuWD13yV7vakyz9QUeIB96QbYt5udJvRXfo28bngI
uywXEgujyPojjCXac0b0i7khwEa51jBoFAaLJle1xh1hPwaHvMF+cPi+Yh2YlYqV
n74dUD+SaumwNzBvsccGfJMEz2Mu5LYxuBifM419iMQNmagfz/LmpOaLTMgejZMg
6EALTtgpz2XxemWsHgn0B1z7Lo/CTEQjctpAAdiuXmQjs+kWiO7AB43YJkIw6IEE
Qot5+74fXovtpBnS/wmJZSQv556BDX/SJDr0kbrIeAwTCzPw9jEYJQh6BF81Z7L8
KlKnSA/RU6urPatsOWnyQMTxf1FRwdPPr4bMNbDbZ4ku1EGu5OSZ6SuGqR18MaJA
uS8g9zW5nx2ZOLBkRpku0i+0h1BRiJkQc4X2KAIy3b0JETXn1uL7rJ7SRx5nHZRP
Mb8VT4At9wWtVm1RCdjuloayCKFCcw/JeJ3TahhBAtjOU88698iqUkQlQOSI/uRC
YgJYiFiYIbX/CGRgGl+iKWjn99xXwWeDzav96us+pnafirrrPvcXgsmnJpOz56Cx
wQmpl6Z5rvx3xGiCLV3bRf4Xl4RojDDDq0AynoX7viB/2dNOPlgAP/daVCzfZQNA
z0e9uOPiXEIMbK1fQpjuV5hnP48WA9tyJ9AGRcf+aeqCZvPnGVOhm11TwaL3oSon
vlkD/UHQW9PlM+cnBHlC7L0LU/ZZcVxpSR99sm2jDIxav5KjEZJMdpTb0NltRtCT
V/sK0Eol/5uXvBJbvSM3uOdW1gQeRUjvZ0rDpqGGVp6wCmHO0mUOo0ZtiAYAdq4J
uXx3ifIz2p5zVBGJmSbMbXb3QrYwduHeKTJt7KVL7CiWF36dsIsTE9nQkrrdWfUB
5HENpGFNzJoqVZvY5u0K6upegZJW/dAw3ACgbeU8MmAMIuguAHft6UDmvwEzgEUJ
TIYCXGmQ2IcoFdRk2lUuP3W85WuONYExWMzcIeOfaxoJHkARaKCl1qyRe21R+WxB
RRuzA8HyJUfHKbgqJOPv/obIY+xGTVtNdzs6k+C4gyHQnft8WHTzLph9GNeEhTfm
87LY/55Gs/y6e+ehXtAMEHW8AcJa5EGJjEbLwf9yKMiK2AJoXSBRHe5qofciBdqk
PTfu/DBi4JXCHJxc+0hFifdLYmXWZm1tWV0m4jRV4AWvpZTty3KD3nMQZgb2gycC
JOAYbtIU2Sxob1ezLvSzzL5+W+YzHPHj9BtaEiAoBtchpFjANKIPtb0CENKsu2ub
X2jjBQePTDMAIftPMfKKRtGDelC3wcs8SKjuNDbDUIbFqs7jRjCBA09X9HTQ211Z
CdkV3HgR/5PaVPCZAd0l1wcxQlz3b55coTcpyGitZUqMy119QU9ducmnGip1Uesk
WxSxD8hX9b4/hYVxtpy3DhnSejkeWgWOytSm6sWLhsPGZezMp2vbNxVtGUkR3rAo
ioZbnHP0e6h+ISfISyCcfYiivB4n7z1+tUwceJX9qv/bwPUrrrPZhNL77//UZf42
iEh12G3uDDZ7+2fsDhiud5cKSNYRRKfOFRLmDXscY4vV6jBHpxfPM1dB8NA67eM+
9FTLUmUaLRdKt1QDxCsyIFGsKW+Lri7xSkBhsVtQQsBo8ptH23zU3ELG2tKmiNgQ
IXuocmc7V2LQGH+oVxAiSvmPaFlXGt8QRy+IF2/wo2JfB8XwnIfxMJirBZZsWmrL
4a0/iG3Be7vSxdr2GRHngqaTxswebMcE1aizUnppX/PaS1B0btYfA/xBdobc64j+
8d/Bciph4V+TFwr3EVqDMO2CPo0iD4yovbvRKQyTvWlKI3aSIQwju2crZuTZvuhT
Mnxzoqj1xNzIlJWRXgYf3vJS0gE9zEJS37sj66giWEAE/RU3ixSMitzbHE3ZH73l
iIZcxFMqC18yI5Js12VH8pgcD5vBWfzLItpXZphSLlN7QOZAncKmOjbPTmssmhJx
m/d2NkIYvNwqjhK7JllCcWq5NgnGKfq3Ow+5761p/5jPpaFrDCMJNeUJodp3+S5d
AM0sP1GjyRRt4PaqWfz0bpF6A5frBhHbdNAPYm5d1PjTiQ8wQdtZvJg3s5nHzBli
wWHNULR4hrNZ8NxHxmSZByA6H8V8A76p9XwnWXSPqs5W1qOXqZQVoGsmU5t2yEKD
evHfWmq8zGntuV3TO599YtrPXAoy+EPB4/rVIh89kGFUrnL+CJiGCyyYOAHRnCaV
LME70WcBdTB6Z3wNHO7cgWNNyEVthHICzKDtpuwUHg+FE+ulWsaM6zHTiRhzNz4F
+vqNnyyIQB5MG43P3P/46qK/e8M0c28Zin8wNSpRWLp6v8MYrG+MHhVNT4qxry5C
ies7/kSmDjMZVpTo0A2/GTZ1hlyf05YY3o7UdZLjOVkU/zYnAorryvoUEUKPmIOt
W10NhlebfEoFe0dHjfAoAEJ/HVi/N6/C738MSZU+chOJmAUN/9Q4LXU50l/2WgiB
+YOT4RdP7nlilLC/b5gm1A066tdwYDF++0/j5yT5kImTqUCLXjPCzDzbvhgsFJE1
NJPaOym4eAIAl6OqyYTVNoLzEncpQDwB6ISetJlLN/680DxINqUyiYQXh7VFhLk4
EW54KC+RbwOwj1b7fp/uuXn5E91i4CNncnOVI+lAP2+m4AYqp9yxMoSPHgMubxvB
dy6qRITetOS9+poEyUogrpb3lgag2OjgEfRt9NjzxCBWcU82yTVAJZ5VjgtmImux
tb2z1AqFL3OExnd1UGTcXfYdObQg7J25Qx2G/ue1mD2S7EGq/o1cxqB6M1te7rlR
om7blaKI63YjZWF/xxzWphVCAbd/8OGq2npa36sYT8BxnIkDg0hb0ACii5XyC01g
YX+sgaiIywhoaSPZ32f7DA34qxxdhr1PyC3NjVuSNgxqPjCMa1OGypAxXS6GQTuo
sq27OZHSfSnkvNb8WMRbWhvWrhn8/a361uslkGHQDGJBEwlBXIunkqsmckHcyaw/
tdCu4V+0kE5PCNryCt7WMTMQUb+cSwOGanjn3BgWLh7GUsDrFjdVdKshnVZl5wRB
oDOsUMF98WP4MHc1QzRfXj4avDrC2FaVcvptJGipi/IiiounYhNkMODD3vZs+sug
883LfPu0DjuTT4Js7/g68dik/RcXBV8p7uL2dp2PDZESEnZhc1GDlpYoCtGZNOej
6bmTFOy4ecunGPFWHobIr/l7+lFmfKrlQqdX/8DpMjyo1dbGtK6XaF8TNqzR0AJd
vQn3yWfNqymBIw4q2HfHpOkcBDex5ESlTQZPbPsdsWJYrDFFJx7HHWaMiUPZ6KZP
bVBn1HOuNP2YA8VTYpGkxplJzMPmOU0YDldvcrBW1loiyN7JW3xqZRsQa78RRinw
XsJ/Awt/ujfL6fCdg42k/i1dLUfpitdwoWzuEgoOoAR8Nrjquadas6pYjCy8hyKm
rumub6wMW5wbfiqhxPV9JVyMZJrKx2NbObmM7JyUlgquaNyEfS4/9/aQwS+Cor6S
kVjgBUB5JZ/cCgMHdL400gKkOX2K58usRNlF3vFCcprC7qa6uo3RqCWtZNRK6Xa8
Ivq+flW+FkLo8izd2NBKRseSQekpMBpo665b9PKaEUxCYtbX9osqeRCeMO8VaPoM
YdCO0G74rCOEH46LA5ZGeKJlX1yXxc9mQq3jEyoK3GT8oa/rJAcWLaLyMvpoM81V
iPmk2i9kN5oZ+2hsEjpu1vqWiq2ZmmSeOtQ04BfknnAUJDnGsY2LQhd7Mz3G6FA2
ppHiIvevOxZhA3znVFueODZlvBMlAcnTAZ5yWdvgQOWSB7zPQJh3ZDqcnFyVoO5h
DUrtwp30h3GJq4xqrN8x9mGKDZc5TFmj3kKkMtWpZ7JYkaezLCVNjVXgmi1lAK9n
tdIN2g5Ap96k6b37WHJOzR1VC/ITL70HVvtPgk6QEg1nWN7P/B0RHxqa7RJK8H4Q
8gC8BQetjKlBQU+mCXc0Oz1kxKNG9Ul4zql9Z/xDTdMO604PGpLqBOfXm36Typ5a
8RBIf8rZcNJifKuI7QPeisdo9UzI9qGtIfxUfToiJ6i2dFuCsawhmNxkxNqXrK8e
yRoCzINAoSXV1mKa+jgnCDBBUqJrzYg90GzgQnAr056wJtC5W/A4lyQ7uPnmhUj4
vX+0Yg6gTgSAtbMu/VoqWtctgnPhV0HWh1kyIE8mlnHamJY5YZflVfXv5tTYN037
1MlPFf/kSueSL8NLT+Qrx/JnKyH2W1kpRvlYKgZqGkOy1E8UFXHKv6x/3fTHmtHl
V1iDRpUM2wV6qKzGSEtogW/dIIqDKW1iFTDyxTayxtmmvEhOFlAsygX3n6JFpVdi
VhAloiDewKYinMdiyFVVErngGlIDt4Ay9/Je2XHNfEAFlSWYjM6VR6LvN0fet7Af
AieMf9GSiNFkOTBuJnXAkmOK+sbhIHVtO3g6p6s59rRo9NkV6hI7RwIRv66B0ZWb
2YyOILKR0b4UVBUzLM0k7Vd5vuXCsNfP5m5uKfoHtbzsB32puYQduM/+vzuiln7a
u9tAPgsN9T67gIDLawytsT0aGyq6Q1CGLvL8IXYIMlNJiJRLLXopBgVQD9vBmROx
WL0QyZtUY6m3Hq1ROxy98oACtAy+N7d66iWw/1bl8RVFqqwT3VVUMdOtRtBU8fUR
9hEf7l8w3bT5XXLDplFh3GkscAMzhoFHdZUzV1BftZhru1fKWW1ywNfzVcpwtdR5
07Q7DFg2P+NXn/S0HyI7BmVZ9Nlzcof0e6gqUHOLz27Uhf2l9ddzp0lo3WpjOGkM
Su3aFyW+lKwa+RMx30q8akyqXrg10lQ+etE2P2W9gt8hbH53ON0d/ul5ZeNxF8Op
Mo7xWvu0tRQNveb1SDPRlD2Sf5tzd3oLfWiENh/xw5fipO0xHMPDch/3jh5dhhZE
ykwReSNdIES1mpps8NABBLce1MjXR8g2hyot/pY741usRfD2M6keN7QFD01U1vJ0
rzUDqnC4AS2pcywL+t4YWhw4HhpBvQGob6oK1s1NYWKWttFdVGWfTocxCkPVdTPU
KSUsu8kD6irJ2ARY2cpnfySjO23Fpw0wS+zcJFaNspHhhpn0a2uT3S/GvHK4gTMh
yxdiXWsDmuSbIc0DRTYEPORkj+irUVNV1k+VbaPPnMeO0KOcKCaTmVezgyYYO9uB
yB90TweIzj60G/a4l0QCEQcOP7T7Zc1olaZUK100l1TsRg3ouSPGIGt89/1ARjlt
1Mvf+K/6UhK6xGdMEZbGugbBPkGMwlJZ8Fe8ZOZlhtrc+gzrhuj/498tT3aCw9A6
vgf21YI5G8lIEZVVP408XZwl4LHRKE1qOWMHMtoegMLy519w2ymv7BZe/n8W0H3K
wuqOQHJef1IkIeFqJHyy/eAj04FHm2+hhkbQm+ASyJQF964rLfNpAO2sy1qb49TQ
RRDTPV0pxjgeRJ4k+puTjopR4o1NMFuD2iflQ5OFow70gqWCvmOQQ/qpkgwZGIqu
yaC76BJ1SkkwNftPIl4n0aZdhGmKgREijnkSAL9mtL7HAs2038fpAfvd/aZ6gzRq
6akaD4AkDDv4rYIWq6P6doxv8KvNWg8DqtvpOLC9UsassuIwE6ING8hNjKrSeO9c
4SOrqr3GWT3LpdGUagJ3z6b6b7Zjk4XVryguZZBe6ah5kzLKKtLXlqdFS+ICANUd
8UzoGZqbxtZ9CNy05BX2ki7vduaHlMGqOEmvMdVtWBgZtyI1hqkqJBC1qhI7DgN2
sQ58QHLbujUX64O5vF3fqDaS+DM/nRLA5Rf2+1zCYaBbnRO8Xp0/Vl4ZSm5em0Ku
hZH/a0aOGxAH8gIi4Ufa6zp4PhAtOqlOE1o3IBVtpBd8FFWSMc34nI2LZbiB7FFI
giZS63hRGL4zdG46gXPe4WDTDCgvLelcetcaNk3A1TXo5Nadu5ILPbw2iH/tt8ZF
BetEp13y+/ZKRRJBNkIadiK5Bsv9EnKAIIadA8ygOY6G2qUuuWDHNtLbY7BP2DQ4
ZkWS+0PlG3DWhM9+mwLboT5cIKbu271yAsM1jq52hzykNJXZNWMZMOM4J61x9I2u
0vmpLUpNWdjbp9rR1P9p1hepmvgtOViWTj83TWUtKCZhdZmhS8dYGUdsWk4ghTDt
pESTNSYz/pwGk1qq5nTRMeiCk2jVj+qMFxgZE6WEMunyhys2667z1EIAQXfe0zpj
fAzKr25dyUEWtfXeh4eRnCtkngyDm1uAZyQyth+vdz0J26mMJB36itR1rMv6Vh+o
G+COpIGCTLfJc+4snmCnsYW3O+b8lJBdN1Us631bVmFrCMyPukqIOgHWw8nP8+0K
fm56ecC81P0iz0EVlN5Qa2xH/5PY8JuYW6HCqKJIq8s0MlQiK1DbE+ssbYjR5qgO
Ur/mJWTSuJk0ZHN57FGoG279U3tg9p/1hsW2w8i8rKUyPrn+/sXWMaR5fJL0kmI4
r1PaaCxsMP6Mmbi1kdxBy8WzYTDz3mfeFLpAU+edTfXNiVL2fpAFE9ZClD2p4OUn
pZnyzjF6eK0Ch61Okiv2uLi7qeiQhoUoww3P3or/VgmA3Pm8xR3KN5ruwM7JitJy
fsgHFB/+dC6RNaM5bkDo8b5QXIg4YRDrCwdW0rrs8ygpenfvr6YnPDxR1kvqNg7S
StCPi6N0H1hP/IQIRNp3tZP+alfmS292QOk8wQpwBbpKRtLtfOwfxMPZjROuM6KE
qs0d2NWRN1sNkyKPOvhYQvnhKjhmYd6/3tg9EoNGYsix+JWKkDFLXPv9lDGqsDaY
PR21vrOaptIngAGj5op8HYcljeu12IbE8hsifKZz+kQF5keTCE+CRU/7zBzGMg/e
jjGNeraSxKJ8fKZXy4KcBpqNfcyj3MgULLLA6HsTU3ocHpwTwrB3vJhNjlvMRVIG
6kPyxIk5ydwyCzdvuL3aYDS3HB+XkySrUqkPlmmxqRMHbD1LCkfznGujw4NR6JgS
A0MjK1RyUd+6ELD/nbK7KRehyeiAaiZ/kEFTcED3IVhr7vbOXbLv5QSwjWMgDt2d
vu2UGEorHU9k3VV6zrQfY7vhpRTENSFjfrOAjQVR7LdW966OUS2w62RYf6ztCsvp
tSTvMgwOtpqVvhn35WnGXBX5eYCCucLb2Xfk1SFoahrVKmsb2rvpoy178CYdGl1Y
ApzdI7v7CLWmneC/eBO+m+E1eRwmR0qJLjBlWOQ7FG+YRrszX0RXUbzOGYFYJq6L
kQyPFvo6l2vDT8GqQlwuF2y6I2b8Hiuf9FalRzbIocYkwLnM5n5HgAhSDkZd7QwC
KpYvWDNdulT1zLog2D1LGoxPq2/F0i9PRmcNB2Fd6svxhvlCo+6DvNSTA2ANJBnJ
cDU6/HhcJ9fGoxpVjsOTDjahZRIIHqn/bef1vCUlw4tB0cm4x8A9bp5dGz/s0f6R
CTxTWlCiBxNMJX/IPYBFXRN6ytGHN71x1O6DTP5cvQO0jHKbALwpsz/SQvI+m9Mi
dgsbUeuI3F4nbLaKSIUhGZekwaLwUeFCClc/ATpU8Dtk82mc8NcYndoThNLl2+PX
vArKgA3DohcZCX4i+PkqAMDHqfEo2dH0SozJ++UorIAuFCciOXXPQtoDdt4Mj7vz
yq5Fayky5jCXFxU0ar6XjXh++S67Vpzi8sKhcgZ5N6xHJ3nOxN882326cUXJoAm2
XE7UHrIrq128YsbW+7uywuHGWoTnHWNur9MALIxGoINKe/LSsmmdglySSe4EbwtD
9URi1kSeJONg4pPIjaaM6A==
`pragma protect end_protected
