// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:53 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PElPmgM9+PW9FO8DVEkLqm5H3paZDOeynz71foHgCw4jXbD2439l3lbYRL5wsfrp
E/K+gZw4rngWBBYvtXALJN3xd70dSskotVeDoMXEeLyb6l552jql5ctXSqTRSfdb
MZBq74K3e5vw59vukjSqu2fVOYPRhfJ9SNAxOBkDxcI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9456)
VYaEZHsTFHFB2ApdbFwc9Z+D4p23bh8f2LZQpidq2lqEKcMh/6OerHWU+R0hIW2+
CVnCxkyn8XQRAwuN1Rj4sLf4Oh2y8WedPK0pWDiNjhjuVWmF4T19JLQR3/pn3MWv
5fdybIkL0BbV5I6hHWcuOxPWC6jaHoamlpteO6mLSqJ4XT5KVV0yJvb5qNNyI7kU
R5Be0/5eWw9SI+2IU31BUkQHHOrJw1CGStc1rHWmYDyjdvnFdxaD6MbNQXQqyjZn
MBfv/niCtdIFENAqQLDuAjJyN1LBw8M42uUCdSXHZDNSzmSO0BPW36pPm6SCGOX5
wFIbeev1xwtu4wDTwUgpmQ/dw1oVCRWRgYasNAc5PDaVS0MDVYtpegwC58gl0agB
J8trSiiL04B2xv/XKv8gTAUS0kQIQYqhXeFe6Be8z3BbeXtQgWRcPT8vgyxH9fdT
zjij+UgEzwebAkE0hRzSJZuxJQtv7qWC5z4kJ994QC0mwrbCdvsJsRoSFSkY3Q0d
uytpO12AJJAyuCeb4szPz929t4fuLtA3mflIYRJ7Rv7jcOwqchodfy31+wNqCDqZ
nOXFxHGnXz1MVW5omeaxpOfsxAA7Gr0UbtY9Z1HiEd0lw1dQ2K1ScF8FuezVD3np
0mNDYRGTFPyLIQyEUTMWQN2D1HSD959ug2Nw5ciaOefSgpCAhy4wOXjO8uKuzjZA
7W0Yw2dGFzPY5tLzUP2lNtSZoFJtX7rADOZ78pxh0NkkhM5HRzwF/RswSYGw0zSH
tGEEdjdCkjtnNxubeZ1RlSS4Y/i5GMXITeOeNUSU0H2/0wVHdvjd4NXqk1KxYE67
wrYI0uOtr/12/hbB5jDsDzv1sKsm9y0VFUwDISfvp2YUtPHv79MVKPs8ONvVnXuQ
AhZQ1NwXrulTS99+A/7NOp9//VxeCxeDQFoNdMpSgPfvrr8Y47k+mC6XArRf1HUa
xJUZP+8pz0RsrEw2j8lJoi68TxLvou8Xu8ckmAEY9u/v2HRLqWzX6ZWbqbxsPR6B
5970ewkeGMiA8rj+pXZrT5XeAJuTFqJDJoJxXWUn7AQj2/xalXvDuEScP0Y6FoOV
T6m25JYy2M7+RQVPKkATsMQsnOcBK+bFoCy9CIXTvBNyCIwnoGPcbpalEk8ILD/q
PwpLgKtOz1msG0qN11UdnWw17ZkBF1e6DPEx0+h1ud+XKaCntvN5UFJJFdK+mjCp
2XXkf5LMtXtj3nSq4L2FspP++rAQcUyhH6AkEPcmDK7jpfMrAeXPf+4y8YU1Ct7J
JwvgoUFWAK1CQ0B0HvGR1DWeVT+9WOutV1MZwt9kEzsyctq712mjsNt8UqmpkTxY
tR5ZUiBsSDgba/7Pj/1V29nY0vtWCdtYeitjppx0/Kmtpjs8nXkLt+ctmlpVmbHQ
Ar7sT928HG0GRG5yBZErM2DvJ3zWgPb5/YoOMwX+thwQE0Bu+6v74BQ+rSF3xpm7
xMI96itIp9KGS6vPe+9jtm8lrYbg+b4NrAvqXPAnwfYyHAMnNqEM/NVi5mD/Cm1+
WaEoHAlnez1aJ1LBo+WMF7AhSHSFQ2Q8x7prFJKi8yUd75U/FqX1Bp5ohR/qd6NU
L5D8hDygzrCXkI+CaifUqiUkHc4I5LEtEXaef37PP8zJFWloze85bAm5Po1LBjso
uC7ifGL6ixkWZsogypl+5OmEF4f6OdRqH8mtUK41ZCBXu50deSVlvRUmLwYdR8ne
LhxFge/tvISk2JmA0uzNnqnLncL3eH0dgYDRNkrAJCGvUyXa9hnpNHUckaNjMcbR
KHLtt1XejraEel14Yvmk0f/2IE5LRKbs0YhusGwf0TkOOy39Xo097RuTxY4lN+fR
Atma8Flq9kjltKLyhagT2CVqH2ulXz9KcP1oo5pu2ZLGyk6t5wQsal6tu+QTCoSb
GZMPDosJ7+z4DJ4Y0vL4Uh3vl2+lMFM0xCdYtR7IdaUPWaXi3gylg3JGYBcKObFP
FNA6JjV+TQ/MzX4F4UqFXuukB7O6tZUP8aXpGdFoJOO2MUDyHMezVi/QD/QXcvyO
Jm+ai7fYlPFIXDbGZYuhoIKg364kXOtPIGQaXvNsxDMCi9sGGfyyUAxVHVRrPyxm
aKY50CtOVGTW31vNhRNqZEyiCOKlsL/SEEZOHuH1Vyotf2/V+2IwSHPE5dC6fu4s
B7iAQCe1PzMa7xYj8HZ7y/Wq0VMHrqDZ45/sOkqXT5TSK0xcuFDCrUXrDZTIGfv/
AzG9x7OgpXCF1ZjAk+u3JZYN2TEPpBX6jZSVAjckBWjYavX8uXZmGB1ScRt2QsnQ
qG9RFbmzWcpjMEFgq8vqOQblSMG0Wbv2pc0C/mXRO4iNTqQQo3g52HT1gFcJq421
2RgOE/3SBqwH3xZmzMKcMp+Up0ahhi7yr1v/WJj8/VICyinmad07r3zzTfj+hsZC
BVsbRTyX0rWu/dtBtGEIONnHkuikkwnfOlq4IW1/3gnTdcUt7Ly2NHRpErZWFTLb
lQ8BoF1BL9I0b/vwtUe1fQ7mEhwyLqiQTXLrzIJGZksfZFkwf2A1tbUJRaoBZagm
KmxvC/2bQyLswZ+44tORvfmVH1tVGzj+I0HFvjGQYw5Y9jbyk1/2cURpIXn9Durj
mEqOa/+ZSwHnH+BXGUdMXuVPOT5Ur68PwyH1QpIPgp+Gj5mtorusDMBAtt5+40iQ
TRKgPQyq/jdsPEWF4Q58gJEaxzyGyK6UxB3/xfbaZzwrCVGwHMQTsNt6YESDuiZQ
hzqFuvTp3FqqizSArmFW4otN5slOycl4y9+jjFuOPvw1M69EtVhC2H/Yd7l0+Q7U
oHa7qSoj4KgTI1ii4LlIOI8uxOORTuEgv74dbKH81kgzUxDjkfqNhXEmWYjViWFw
8Y82pUKu3JtbUwrti/AYWk8OJargOXjUv5unCKChDrAvO0UUlS1h5GVaoDPzk1F7
gmcSiosabpKbzTxSOJR0k8lPDUff6hFPESYD2SAKTuoYFbCTFWev9mZDJEgGtxBE
VPgM35iKT+QEzOhk9co/ZfFSEABnxG9TepCNpiz/n5HXkpv1MTiVVpx7bfqTzRBa
LCyDdgdvdiqMu3wmEjjnMHGcvmHzhE2ni6uHTfxReoiTE6gl45RQCMWU2MSIe/Te
eZZdg9HSJh/PrqrJ0tf4yVO5q9fidzWagLzupgAoHd4my4UtBv0fJMHXCdifCjuC
cCizaUegDeUPRxC59morce7sWvSVThAxYlpkj3ifXN7cqq/QBkjbVq4rNg3PQgVY
PQZkiTix62pvq9LOE+Z4r+ppdAf5xR1rTgpYDCSjLIHaX/C7k4hXKVHyR7lgZ31V
qXnKt3KfgxPVkSN0JEKnfLXv4xyC+a3upN1gfq3v3vDHeeCF9V8rz4LK8c8YOQKg
H5NAqMnEilwIY5e5HdZK8f+4mlh88T/3Ogv/4t7bJ3/1tFwLG8EfR5DtUsKHZuLd
2B4iccTo/3K4SuHUdiqV4rT0rxA2lVRbKe5KwRx+D9oWj0PUHJ5ZefKgBYFhxQKk
vBEdcFssn3FizvbeiFeaMsJKjs0rUlGV4s0INTaNcOhyyXkO386ZNxhhN8wRofUD
DezOafEzbOA45+fAzlUugD2T+Csz6d6PgS7ACNpaMzxMV5fGzJVlUtX8nXmMy3Hf
/byPXayflS09hoaeJ2LgDe51kaX2ilxpHLxs0sE7nJVYRyjcieb22TV2uJ7naDOk
+sBIteeFlCSen9D4GFXNwksQCcJTDAh1yVhqSPFwrJKLNLT83OCbday7haJGWdWi
EhL+pem4uVLHA9UICwfjWScW7IwslyCIqDWcr/783IBsB9BIzQvr7SdlfwpxQzIJ
eBDjnyScDNCg7Hw4nbdOIAtLePNWHMqc4z13bm96hOEqueKrUvF/XFA+yBFZFdYL
MIdUg2IElqtLbI/PBAnHsGLveifnQC62MJv0Yv60uBx2sUZhzSL9lztG0QVZYTDi
R+eDG6+OiMw8gcNOIxo0OLJ2WBSyiWiXCZR6z+gvUSZZjSnDZ1KeanqEauOX2Lyq
aUSEU5ge8ae2PiB+RnJiePdJojOLiydd375ck1FOqi7wUcalcgu5BgqyN611I3OQ
xQSKP+obOxTj7XKk6wmCB3B7iuyyEc7qdU463WilU02XepQJshWZeUfzz5CbhLUr
6voXDkn53JFvWLVFWK+DYH8YjwM+8Zel7bq0erUSccMHgwH65kAcp3r7fzhek2hf
lXWTt+jXBR/zzI7Bme3O202IzcYlKpbw5gmb87wGD8gteY36j8w83qqXfi2fQThW
HFostjCQloQqGnw4RMnHe1M7X7pTYmJFANxl1C70xI8RdPUh0Kpj26gHPOHU5/OE
68MKLNdHqGWp0WP+n607Unni0cNupXpwXULPRIEF+55iL0yAqmJFnLDiGds0gK2y
juBBhCGnC/mRc2V5cOo0G21jIBQjcLy7MitVE7uq7J443wmBJiy8rSrHlopnNkiQ
ms8jpTKE0vGI6/g18VWfx8QI8QQ5iCocDj/Iz1ittp6h0aogQcjRoUBOGduG/+EZ
3lgm8otXn6nJyrk09IRy3cOV4F5JpXXLQqeUvNvvkKgEsEbe21DGPSi5/mUgxQKk
Kr8n30CNx26zArsQPvY0MLAA6aSRVa7hGhnNqmHglGBhVWj2myOz517m+vRmweWq
TbmkSep6q1ioGuR311tNh8Qh9JyZbU8gcTQpjLsGOjnEw0SHukXozBtjFKsIIz7B
N2xIAjoB3nRGOmnBsRDWOEyA30IsCbKlsQudpngHyhwhRXaupQWYbkl9CJgnM51q
3VDhjSAJwcs115UOpS2oPc2ei8koPNWF6F+7uE/wQJSZ2mwDUBf/jls6q16GgKcF
iJtUzc/KdpENqLgW31Sb/9MoQW0jYxD5SHgpM+QyCPTkO2t0VFNTMdFzmcemgppv
1B9Ua8YC2iZx/TNGMYskxn5lR1nA7X3//SmYE35A6g8Zm5uS+bzvxTivmGsh5Nnd
BYozctTW1ncqMo3mpbZAcY4gfuVfX2uMzmnGS16gARsBJqdejQHOQw6Y/kj4XVJP
gdRCfutsChiRRJTBgSvEPnqSc0ASW+XxSYgRlR9ubNB7OnSUQtarHMNfDl9sC1Gr
BNNZgZmZqzTdGt2KjeAH+eQVWNBxz2a8uXka5U+4qydkdKffVxhQQnxV1ke/d0FM
r0RXasu8KL8niSps3QX9NV719bTn9uuCrftTJzCjgrpfKy9ylISkx+sbiQYG2+Ox
x7PHNUzs2I5wLqGj83qGtDhclt4b6J2lUSmTqkwATgW6hDag6Nos+vyuaXkHv+V7
T3wYryHvrmMQSA1iQ1e02Ziq+CKScUclj8b3nAI/UPwifK6Qv/Ph5+pKsJg0zyfu
0KwgAEM+Ct9uzLZuHOwY+XKN/zZLDie551Zzx/hs5XIPF559S/ut3qb5cdhdBpx8
4HGcRq27ZSZMuG6cG/GXFjwXMDcTaeBeTb5RB97VCfSi/SJojCBgnRXSsZN/OD0j
i9XTQVLN2uafbDDnFQLbJBHfv06GuMQdfjz7yXLeuqMJmA/9wgCdBVniOsXQnbiV
yilEZrAZPGASLQXXPn/vFmiBHzQj6eF8jwPtduH10eeC4/JCGGIPw5ZHg/BM4DOJ
u6Qhlv2LF0+cAdPn9+fZEmCEXymveJG84Hz08mTxliqmIc7ldbKL73bVHHn1Wkwv
5fTAzKy/uAu/IVO6ap/IULorg9q7H38iSYFAeZh9XpNxOhU5wcAfO98Od6aYtqW1
XpSV+hqr3a5/CD3rSkXWMMrpq/byDoXv5fsJ29+adOrp3kAWd4XdpfTc55VbpCpC
w2pf0f3CamcJKZMs2arD3/7d8DlRKpLQDgcEVBXCUInxTJEt+p9ydgbtB1x/39+r
FVUq0xMCGCO7Z4Du4gM8MwVcXyaBgNjXhaI5NFGClu3njKL6swyCz7chpxnBV/tQ
U0Z+mbDKkaPsG57wJ33do4k9v2NfPxBjqlhYXcpsUqRFAd8kHpFHXrkSkhXgZPu4
/4GOvEWTpv9dqu1fvOfcw8T27AOhfpsigcbRW7ZIE79+IiSIT5gqQ20lJQeGBiT4
WX5dOUNzE9axkEUXOyax55s7/71Lwp8gdrN2pNOD8GRI1tH5kkifIGOuJhTIVZaM
Go/IOVnpIfLXRw2WZYAVVSJbU9Wz5dfVIk3GXZVMANdCcCU70ETXGBK63wHDbfAN
lvFsS3TlLwZ6GAIzAi626mpR0bVO+nI6gATna7LXaszn9tCMwIAibqRz7buR+7b1
hdWOsFP3SwGOCGD6VlDzfWCszoF31SHrnWp1Saj0B29QSGBbWTAuzPJ0HPqMfzfH
PLJW4uL6u1DBAYBvTX9H1DuAAGMoWO+8ZcprxAj73ax6c/4ywYim+iJ0gnRGiZ+D
JUYkPr2IsWi1mrxEHx6O/4IoksSAqWlf+CLDyEPkiGO7NKXu6D3KmnuYwFS1bh5t
hkpw6oMfjmAqsxX613S9A6YmQUxrgfJaD2TwgeTpqEQZ+XxHxNhJBUa5RvX9wf5C
3oRfD5Q/ewPOwFoO8iNREFifCiRfaRwBNI7oLmq1bxQk0Ml/KktNYAFozp/nQeUc
0vA+hBPtROhe2DNIJeAR5AkntQkwgYJfNBaBSkA524dzumBFYKYtohHXQT4Sdh3w
ddVJAG375+ay2C9FBVII6Ba7sfAkqjlfEzdJkVoina7tjLV13E8VI5vPNj7Fcv/c
l8365MpuO+46cMcetofU7OBtM/d4yiMiLXD6kN5VWX279Yo6okTwpSIQi3IohT/e
eW5cbC1O5SCII15lKJ/EavCtE8cW1+GuUv4DsBsem41vRZq1jOKSdfvuDKTRq7kb
HqlDF1DwylIcBhS2/BLVFWYVBqo3KC1QoNozb/IUfRLjB+Lu4Cu+M1RgUPaEbld/
eawN8bWst1imYOiZcIwV/xoVjYmpHc4Enl1W7e09tMS1+UPgiIeFeI5HOqR8PtJo
8ci6pybB6QdtroYLxNZkKLUjHGegt+C0tIfxZRMEXxHvE76GcXf0CRwcap+cKsnO
qEsB6MAPmiqYa/FK/HHC/J+/gcEnHi55eR4hbBBPX7k5jVYGNfBG4s+3RAoC0w29
ZlCIsFOYBC13JW08/dv0b4t+B5OW77+ddZYQgfvpi0UT8xHMyIHiU/ty96Tj2VrP
xfHVjbjEvBFbWTQyYUJiOnwKThWpkdvdPHl5fOnNXg1+gd7X11Oopa+Nw7yVrwfD
zFoOqYlQtF17H3YUx5EcS6nzpuURLH6OkOwPB0PdU2jWlXaXH5LQH/4y38j784QZ
Xtvrx0zTHkIsmvYCJ0nxJK1rMjyzZVoij/B37HkR4lYsAY1KQ5i4Q/5BF+U5B84A
U1RTZ6hiXSAYzpgrWjBIr6wEUKXUvvHpGN2snAqHr6ftYkUB6ubnOku25Cyrhl6/
W1bU3u8ZMXF7+cQ4B8ghkY4JtiqSW7C6AJHx3B5ST3HZWlic9cEmRckLdXJPHKMT
sFYau188g/6AZzWm4VtuwgpixwNCkEemxP6SsC21kyvV3shC30+8WrHQT6GjTijg
7zmUgzlYEYqFZc3UdNhtEyr64MpB9T5CL1AW/jSKgdlfwlx2tdootcQgEeTltN/K
/5FcCKwFNxFrzyxxq/kaCnhQVCMmJWTE3S5RE6qmsTmClKmvB+2Fv/HrpB0A7KX+
Ms1hvdzNk2qdge9uLY5c0mBkUZfNB/YWNA3WG2Ge18xr4BnH/67Lha8m9UT3AZrs
DgxaPNnII31A+gQZpteQ8+vfmFv/hFaqsNpXjMdo/nPzdLmXss4I/83MH+cLyEKZ
DpIwS76SyxOH2WJsTMSWrTFW6SlmBJuPfepV3JnU++zsO7g7Igaz6U3uPVAoIXVa
PKmDUJDDVmsPKdYdBRdpKdaJU4h18tIt+qN65IGhl8BTobVaicVIZ63aHPKiid9/
GD6Det4vluwOQ1KtXfOHDAYTOqcKPM5/qAZzkV/XTJ5Q6juDDJH52zNqbWxoFfmw
PkpDq5JW0iw4MhJQ0rfEl27RTuwcMmdWB+yyJaBNiiwQjTyRHEmDJ7vlmzlSFtSb
xOWQzKy6ARfia+/0fSNLs/u6vb8KGtv2mkFs61R+/kKxB7KuT63CdR325e0guTXY
1BvbI2WGSSP4PGgrgCzrs6N3GR+JYIc5uroNUjmwDvxsZWB2s+WA0UmlVeaMALB4
1SxEJwPwnnx9t2815yUMk9ntd7Ergp5/ca15U0+yrHXq1JPC8Kb0pbadupcISGuE
EzphMDesBjprd2ChrJu6qwp//TTeEO32y9GLPvC/flbQvf1+WcDdsgohinJgjtsF
3/PBZhK3LVyeTqnEcjqgObLObtoSE0cf2zd/6TFMChHULPRGbayXkzDiGz+JvBVE
F6Eilo/B0ILhJ+I+wA5KyE1KjP81dmr1Xq6VQb2hL7SFxkQs1Ewkwz/4+U/vsu7b
UOZllhcFX3rTSfWXzy6lv2ZBb5TQi7Q+CLxWz2xHSftfuVY5BKARUmFz6FuAeOK6
FvH8T1vzjP4XgadApkT+bHQZwk7fjRlxsADaIdfOyaHCQRdLmWrfIeVpfL/5DjCh
/g0U/HR6qyh1DMKBMN2sx8MRe8TxpeTGMC9LEKAiW1u3XoulBuE2Ao9gtpgn8AZB
+gWvtJTdslCb6hrD+WfDu9aJjVKfHDDxhyivCzQMkyzWIy7N7ZVAXvKSVdFeP2zF
PzgF3JCwNAdnSuZ8ycpG4HBMsV4mvOWr+2NAUbDT+ivibqF2RVDYoN/EzNuLQGhl
00ILXaMGN+9nWnwKsZ0Ot4byBkO8PYW+p5QwVLuKU7Uvp6RMoElo34jtphK0/D+g
S+4ca2d4EYo+EIMAeHIX7W787ytvcFGDCh5Faf9xPZAYMQkC88Auc/bMtqY0iOgb
j6juBPaHi8AdgTgyOnE1J7ULVNK8ObvwudDOh9ZTQu1Y5UbolgZZjM00zsr7aA0w
xhWSWG8+4Z/WG9K0ytgHDMv8qFt9iaPSZuXaYIr5eVVjDaj4Fl0f3FZSyN9HvxuI
FQv1vQOSku1xbEfneHAG4z/NtBIOsH/eHsLRjYtg0bXoP3U6K7t3rYHAitt3sd/F
Cq0YumMtbcXX0X/cKCyJmMVLGLtPKsa3Be9eMt/VxP9mHrh1BCJdxGVIxsgs7+uR
crLbYbv7/u203yskRa4jx0XlyTIm4IJJs4i0/RPve4ZGVS1dAGa5CORfYrz6QV4H
TZRLXk398WlD2t52ZDk3Yb9fs02UYJNwMGYfqokcu3N8YTK72S4XoRPV56hnwVo5
cYpHDBzJlJ3pcVK9YGbtRoanAUUeA/cf8mxeOn+a5Sh2WhvfnX/VE+3ogM2V2Gwq
JhK4fq25QwKFQA+u5mYdwCSjkXXtItY6ZEtsyuuNYI3Iley55gqr6bSXzFfIsRly
U7wDKniqgt5vtpdDheofmSvSvrcqNdAauv1321XnQTVLyO0N8AgwfomMiAZTWuM5
Ix33dY/T0JT4C5PLPZ6U4LCwdZNJpz1kF1oIOudK7AUwhbImpzcMJXtGSDFC1o+Z
QC692Eudzr6dtKsOWnq0OiF507M6oGA3GVjczHdWndccMmD/eDSBgwFHw2wXzmUL
B48MUBBkWmi2EBrOUeAkPYdbRIS1G+BeObwIKKLnW6v+ZwuBPuvaNfjwEoDXk0rM
c0aFfkyKa7iI1PrHok2PLHUgck3cjNIa2rYHrxV/9LO/5JVY2Ho99KEWNDLeFPo6
ythDr2mCxtNfrcJxgSeKgpdxFrd9gS/9Hw0TCrek4tuzssAzw3MQyBnLlNhEHRDs
pZ7Z28xzlInSaojNXNHMLoXOFx5Y9BJyqoX3oiWJDJxr1D9bnW+qJUo5JBfqfbNC
JOiG0xyXAdmDQj+++LNNOhMZhpG5YsoojDpNjWXJScCjDALG+FOckQgvdIdZ0utB
6WOwXjAROdw7xSRSh1hLyOA9dNZE7Y6g+XCiRWAT6kX8PlVmBjdJBBzIQjNailGq
r/j9RP2wHaEwZSkS0y6oi2QVGlzVmR1wcljQAgPKKBJ6vc40MgSh01Q5T4rt/teI
TqMU54ADMmkNfc0cg9taveEdLV0HguBc1ZHMVp7Ob+OoXSCbSpUQFULx5FUtHWrr
dyhgyuj/pfTmSaRlDlIGxg/DazG6wVJdh7Q/Fh2tYOaGfYuYOyh6OGprjkNDiF4W
16vaU0q5Xg18K0Up/sOH+IhuizXfaK5fTeYd8A6Pk2+aVhdnBQ6nZd4L+1jA+SVo
krpXwBrtcCtQ+N5HRdnX4VVUhgVa+BBSMM5D2TYeX5N3T9mQfqbhQPP7bBZ0hoM+
l8+xFH/YHQfJL8/YDrsaFzmPmANojzQ6H+2t5ijlUSAN3EsmLpcmZQYVu0bBg/yt
rqDF9ybYW6bOiHvO9rBB6AIcXrRNVlhPf3mTT753ujS7jyDBvCdrw/Pcn0F+gQlf
pKFLfTgu1fLTXczT7Iv9iwRhNKE4YcAQ7uV93G3zc3HvpP2+BU+Z3aG6Cm0IpCJT
jVBJd2p3NC8IK6id844Gp58HHI/ZzYpBK7Nk/9MamDpOiQ1ljQ5IKjEgkbQqksdP
teGOosP+NP+33NOKyWPrMeIyjWqcmz2Gm+sbbQQZdJq1ifB6/gSp2r/xj0vLUvCM
kU1lZl77FJRrp6iisxg1lHte3TCQwiUfcjk9rdVq+rWyMcbb5yFchjJP3/RWzUcd
Mi1fYreB8Chtp79RZLnTzVJY/uxfN4H7z5/m1Q+antFWJ/vwlLmpjIkDI0t/AAbt
JwaLMfmDnpyTef78oP17XuqCQnoamBeA1BcsSfQ/wXxiqnCUFG46oma4VZ/vPtfF
ugE59UWmUZzWPpa67R6JYZz+l4L+wot59A3c136b7QrtmsWGpVcn3QlMc7CaAuso
7OdD45FpLy5nnMEmijkotnTZLdyyOLbWywBjpsT0KYgGARaOCdm8VwD4jhYXe7bv
CIY4ClYCQ97v3qT+Bs2V/x8e+WnQF9/gK/bpDlPWpIivi/sHXJ8VuZolGC8FBGXN
VkdSYMtiIykzde0QzcefmjSTdQnJZHZBh8rgHyoiuyaisomFJZspMGjIYW90JVRW
quJxOfH2o1R94pv3v34zBP1rRJWXQbdmKofnZI6pbZFyBuyXJhb2As4CC6ayMzjE
jWDLwm/ys3DjxKxW+yeEShk5BgwN7ONn/tOJElb+17edOb2/fETsG+WsFvT4SKS8
0Xch2IaGpspAnotbAyNtwOelh9zyTYHuVRp73uXFOkg6Tvg3tW5ZDnBhn1v9U5Wh
M6PMEFrE5inu1uGzCgGZr+HsukOXX8AFYrc1u1MwghqqzPVKBrt3+luPwYLipZqn
TZ850AijeCqPZx7LoHr0z2VjKpWGIuVhigwxOwrNsSgffheE8DCmZYCVq8e73luR
05hXzGMSKilawiDtMKhSvoXaAFEoER4FqdYudS4Vht+flZ44vEo/xJCzRHza79gM
Q97YSevu7xkKBrulkHL9sAPojKGQP8urcllzc9SpKDzZZl0ukPbUeKlVCNjOwqx3
5yR0EsCLXhsu/1u+fn93GozuLiMxjKCHMbeI+XwAH7HtviRhKrf6y2zwGUQmTOVY
4aWxmWo7Z/D3ljq/FKwmPEml6G85GbBh8qMRXfolS/NEWWIxKd8ZLLVaM2ftm/Oi
CJbh+cvHDrmUcDBn+m4t5RP9W686etGZgAba0YBaUBVmlLONNYe7Es04iPmjbRdO
xrF70V03yAeqg48+gmvqGk4BIsAjMUtck53sJMCQ4wswFXeWt4ixrV4ryt0Akprq
fIpK8NdsTN2uPYLNWqWwOWmhM1jhu2sDoRGUhADIRdi3lO9z/ZuJta49QnygKo5r
mf1RoKM7eygc3JK2k3lREpQmnYMjDpdVDgAN0ww44injci1WIxin1C6Cm+LdZg7o
sMwOZMlYMTYKQGKbaBwfGBkjsSxARSr3kramW13oNHInd8O2eiSBIspwrHxsUc7W
+m9TqXTTh4Y7DgxeXdh1Np8ZTRJ5y5bG8IWqni2x7iLl4HAc+a0sIIglm5JlR/42
5+shrDkfsGWdW/EoWEwir5MYn5o7ck//CYLOtvYjVxKcWlvt2p65x4/BnRgOvZjP
tIkl8+t3kFN/znTHcyxxF44+zO//cohlXUCFmnluLAY851o92F0rIWpCVPAryPtb
RDjoXUE66eLu1GCU+9n47nKySBnF2FaSZBvswg8EH4B5lwYZV1sic5ZFz7RTvaSK
c3NY/16sskJBvrtuBjLNGtCF/eHBbQn0Kqr7hNnkcY0Noolh5ksFoTu3N/Ct1m5+
genMBK5XzuKuAaBEyL5/GsatQEtGWmH9ltLd0iP2l0dJiHzllwapguiLTMkXQqRT
A7vFWVPjj1nFa5bKEXLuS44DmlzhMDGEvUGyYquWHGjwh9C7aDevLXPF5U+4vJxh
UJ7Hc98ltwfaE1iDJdh3JHr2GFAWlUW2dj9ZWNjE6RXZjhUXhEpqWKkozAMn/HcX
Vj7mTkVeElaP68Be9KrNgpFiWiJpLiziRpTssGs4obDHQLENOVh1c+yb7AoCgH2Q
k5rKbTFFDytA9GnKyWuEyZ9CNJQ1pwcQpUDZ8LhrH+HA2UuujnfyS7oOtnRg00ov
`pragma protect end_protected
