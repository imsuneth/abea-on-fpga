// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:31 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qh/+/UDVeoJyrkrRbIrZkyI3ZzHf4bMa4EJ0qlbI/w4gkMN+BaetSlOW/x35O8eK
TiV/sLuHEn1pVmEojw+CfhXAJPKGFe938+uM4SHcRGveL3F06Cg4mhIg0BmsPfV1
kWUAtgR/JXUyShatiZnAuzLTrc2cypQ4IJ4pkqVhr4s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26016)
lPkLFB+qDHbm6SqbIAjK717/QWGH/7CFyu8SPUGLpu9QoRrQxrNbYrWBEO9BrjDM
oqxCj8IU5mfAiJ1bn6ml0DbG+0tsqXJ0xXhKVakD6x5oqK/5F9w2pcZfkJgQkqXY
71M2djhltJ5avxk+4tmlIn5Uj6CSntJcdboJYPAETNUrycBXICNQs/wwPWdB0w5+
3WZv6G6Vu060J9cFH78MhYniMpUegK4BWoFUj0zG2CyV8HU+635thwzJ4SkAD9kJ
dmVZw4yjezHUnFKnEvr1/t0B6RJAMVATXutWdXj7yrHQMNzCiJipzbJcBQ6AiyL2
EWoAKqD3UpoW/SZOUMxlo2j/Qyba8hLiapp9ahLeo/e1JLQpk/vmw0aVv/khS24X
8Vn5qCrbDfxHcmXV0bn4A1CpGgCnla7zK76UmWbQ6id53TpfDs1+pF2q7jhj9lRV
Iu6ek6SCSC5+QGJ2zQ88U6lYoVvGrKIVLga/o/f+tcYSlPpiO5zCTQMlfEsV4GYw
nDU4Qo4fvTjAzZfBgEc99IyLQcWfjiFY4PlvKEZc8AXm/sI7UInaXZsd1sL9I511
xWPAlP5hsTXiMx45yzyMCYHu6GRuHNyeCZD0byJRgONejzriJ/ZI05t9tqIGg7oF
s7ilreqzpoZRSg0g1MnPwKsks9nFghdEO6J/joFrY45t4czMh7Vs01no9rWZAarh
SjKjE1eRNpFssvEWVZypakrlErAHBIFgodTF7Yvy07uAsnVZkSgP9gA9zEsjrdQv
3pmeYKSZBMa3naccRbigWYF8F682s2sdORg+C/+YJ85Vuk/4YFYy/uEC+62UpM6S
oRgyCMZX6geoioZ0CxNMhoVB7NkukKfCVplJ2BFh3j+pCk7SSJO9Zjcm3c45JZxl
lz2Y4p4pPpwvsTeX2DW/hjKGZUSXQf1q8VB7QDHlt/TLk2I6nXPbQAb8LQ2wDcY8
MUU3Lrwa2yXS08eSkSxloRnPA0iUGeDXHJcixh207MyVXDWPZlvLPTTI6GdRcumT
2KTG/3XDSq5+cyqJofU3gVchUp6psPSVzW+qHHwMQGWFRLDrELiBhE2k6csB6fWS
kXYMzWwjl4Nwp5oZ9SLWKdfng5YPyjxIpSfxjfQYSsVX6juehbCEp8RE44tIQR7o
6yUtxEk6IKAv4OoG6t8uQX9Jwiojru0a5MdkTM1TUg9gXR0Vtf22/n6QVAtmAL9T
SnHC8B4dim5DWCSi4b1IvNZCohLirLtjSdAjt6pUtar/z7j9v3uMvsiF9EwsyUJ5
edMoG0yzugYl8J7c7a9a8kaQWo8QAVIWgPCIGp4V5kHG4LQIh+mitj1mvPSgkXFH
CSLVXmQi16ong6Y4J7GnEctattXfJMXEVLd5l7j42g94NSNmYUTnRhorK6V7UQgd
QB5y8Uuf98G7zJ/YL2YAyjA1OfUyQ6AcGQWbww/9Bs1nnLc5m8d/ryv5GuD51vgq
miFqMlq6AUBL/TAbova/l59Txa2OZ/LkG9gxRSSAg5Tlk8kNcC3iYJnTeL5mqqcK
YTVcAk6rRKTDaYz1jCerffS7tFuAcIjNsJu94LcMsjhJRlFptvWbkLhCupL8QKFF
PfKxdS/D3Fpp05oTOPHtjv1tHYJT6mOUoekk7tVnROooSENl3OmUq7AyMv6wRyiz
AaBPF+TdrpCGeTKMF/oBSwRui4gaQXIV1OkYFF9Y30vqJjCtAniwATtwnsdB5BRG
6ikzmsFMXDM6Dzjfpn+4M/RGkzyzfzB+OkNyojhPXGO45Y1iXYT++3VO7NEoM2Xk
SziBa/9Su2K/AOWnfkCDrIkIGv7P7xj5P6AHRA2VJ+ym+nQpELgJccy9jysfUnwp
zRshwD1jrtJO3H6n6H638t2sASs0jx7Qd489fX7HsbBEAko5vgZW+3m0EWhHwjsc
8/5U1d7PpR1oR7OimgPbHUR4AiYrjx0+IzasRQKxSu8nMIEn/DfbrOFjEUmA3saY
pIn7W60LSzaXC3LZ4BnURJVfY2zAHYPeU4PRfxe50LTqUOTVr4+YSMEbjTE8YU+7
Q0XnqUq2O42xNh1Cdgvz0a8OA8TG/YpJSt5zb2qjVDrzL1m5Y09dSaeW+YTFIfQ1
jzVeOnxvsLlqg/GRiaVJhIZ6gHg+I1wFjtT2eLr/3dmZw/G2YuDDYm3EWICxH9Tj
gGpiID3lDe9S/GqPGNBDj5wZSKSleMuaf9cVnOB/BAvnxdF0VTf2RTosMUrRlCf/
xz0dr4+yqazV8O1fvF03bdRWJnXa/RzQb0JfFa6jI4wZNvlFQ1qfed+6lGRZyDYn
I+4EGqhI4awULu7vFy5IzNSZ510asCmAA+Y2LZQqOcz/XLwvBOadV/XmTLm5K+jV
AAYTXD3fnfrZxrUd7Hf9rxdY3IuMY4HjJV2e/NxhuC5FdXfTaGNW8QyA9QeCfZ2P
/7kLIEFqliuuG09XPGAXHrT780h+BmY9Ziw0Ha0em5sKLU6weWnR6iDi5vVbEYwx
RYNFijSG1usZQ9i/CCklJavJ3ZGb/UyxT7oxAckWDD6yogvfslU22yguGfGqCteY
w+DkzpQZJDQ0P+nIZ8XNYqc1rEtGGpz3yN24SDatpbySqNC6//bk+gGzW5j3QE+1
9bMKusM6IT4f07AOYSubMn82b7k3sblaPuxi3xS6B86UBZR4m9lGczfMGdKUyf6B
BXPOEJp0HO8N7pRbiyy6KffZX0hZPslCvkGqfdby1fPUKqvZi01N+TZrvjoTnmlN
Zc3Td270AXFAJfgsPGaQjUegHXJb2wH1gMuWWEzZdj+LuxA65wNptkjcKj3XiAQB
f3+eKY/oFSlPg87V9H2k0VB16T8ZcMQqYx/sD7fw1oWJXttJo/5pAq2o7exUW/LV
Tx3yb9lI5pha8s6xUgaGz71fZdE+OQAZbEXGhCnltoDONxEXeoGieHXF/64SSqsB
DXhB1w3S3fXVdDgj4JC+El40Jb3T3UFuIUhA3jTkq2BcuAcJlhZWid025xBjuUmO
jQeMBilUzzDtCVOcdk43+MqRwsFQpEl+oy8Y0GrmTi98HS0Ta6AwGnS749K1t9FN
kQ6R+iSSMRBjVhZDAAkLV5qmn7r1+U+hz6I6gNB/ZmpGE/YYBRYPq/F3FWlKw+3/
YgC2KrlUmli6NTfG5iTWsHTnRSXE2Sz4z8Gt9Sx2+LJZd0oTnAnQhuKcW8zBmKCO
UsePR+vfUFEXjoJ3R+75sHq89FdSYzKE7SrgKszkqqsvFSwYrasQPEDWMFk9msEv
MRgNT6V7RJWhIqaRQ5nSHVwlUUcthg4yS3M2VQCrnUiKgh7qn8+NldRhXwgbmLxS
ISB+QVzOeci1KybZ5fQaQ3c/ojshYy92RCUL9QMGGTciUNieARCj+7y3ZQ+KoxZA
dwue7RC92hn1Uh9HYaEwsbd80OIjguDT797hVWwgklRhzZWy47F18EtHbDqXCIoa
dxLmaUVz7HP/KeU4HERRBvD/SgT4ku6SlLV7+9nWLnjq8Ne9C8E/FIcq3Rj78AZz
utKY/BSiCx7v7f5aguvrZE7lzSuKRAcxaBGKKGVPa3/Mtz7pPOApN+F+wWH8PDtP
HzmFmum3lA8qCZ/5urp5IDEgszibS9VixlTyi5M++u/vcn3xGk6xQpjXxPPjBe9m
AcFLSs+GQqOCjN1ZHokC15pAGDZ7WNrgiJr7B4AUuFlPWt2EJnGsHbKf+0hNjcTU
VhxXESBbs7O0c0XiACdUTW3YbCx1ZCD/6xcowCG7iKCG17MKRqf1FLOxXTaGya/1
qsc1K4sOutFFwIYeC7zl7E5DTZRZLcVtSzXdbrfYrJJBkOrEO1uRB2Z83npfadSH
GU/3YK5QwEcMntnuE/Z05Si1j53Hm9+0bG+u+NXG3AVO8KTLaRAoRq7PtyT/Dlgp
BQ9cXaVyHIVOpNeFVwvGhzP96HZfzhOx8fGZMZUQbXJxjIkUdIALNf39pcFLhrZQ
ujfd25wuewn65SQSrxT56Sv0h6iA2tgOWoDaIM15aZk8D4ASg9AjmIjW1yWLPye1
G+dxgdcF5d7slqgnVk319OgiYD/X03ciw9vxLXIC6PfMayw1Uw3dhX5PqmaMKvRk
rBkK0bii7bXJCnNGstxv7I3IUwXe8QeQJO+ASL5YWkj+6yPyag8dRrPnYcTfD3Y8
ANp3HycZlUIHscmBApqrlJ9CO8RNFDmcQyPGXCd+UdajZD0RBQ1B78lAA1rhsa5Q
cI2OAX/BYZP6kOGlFxKMQ8rJVyMS84Q/GQmaQizYbFl/Ft8xeP9aaSmy+B5Gz+HX
1U21afmF6tocjFqCg8hg9vZu/VwMzvcCFzwZmQDQnPpFlR8+aqGSKXRs1Xsji1J3
kQSBCeDa4u/mg+qXanev03S5KX61nDkEZBSVDaXXFx+q8WDHOlo3N1yJ40ptfobQ
1xhQLQMJaftC/5v/zttYuK49SjpG7+dHz+mIffHgBL8lYzKitTIOd/k5n+GzYraU
WXI/rroWtUGN+MANjxtjqG7aTVPDSXFaoa7G72l+zdOPu3U37DWt7/6sx1dxiBGh
sFufHYDtrbocMDtVI5139wg48+36yGfZvzLmSD0ngoIWldNV3byyL00uDH05hBQf
KKPoIE5uRm4URUAvV3Fbs4no8ZPxLnKh8Kj/hNPXVzFei1DJqNfhAZyfBH0PRI1n
xbfy6tj2El/X4W8I6ThAbWdg65citmDdHjUnHA/N8XUHM3T7L4XFI03cnJkahm6P
Iav3AU4hA4KIuHp+eoh57fn4971Om1RVmOMirQLp6B+MzHPAQaaiL7id+u+8xa2y
PdrCKKqUujNcvOvr1sGgN0U0Kae7rZ6PX6a4DoZa4JCYypvypuivON/dp7/TrQN4
tzd2L0jW4ehvgFS9tWwBiDVnDZKrAWS6pgyHmcrjW81xNz73aaYT8wx1b85zPqEt
aY0c6MlWMcNyk9AjCjAc+UGcbNMq3hK/6xlTr3up7lwzbIZ+Fu2Dgp3EhUvEDAQc
sJ4uCKktGqGo3gDXl9qlOjJcW0kiXIvXUTOhB1pzv2FQW7xw718gTyFu1EdIkOgd
EkE3mfMMjXLMG2p+ptq2ru+vVopxV1RBbELdr1TFU5M4DwugHeb1mhaQxVroJI7X
Kcuu4os5iwEgo6OfbcXMbhdgyRP9wnqJV740ZP5XzF7Ops87Me46f0Ykl4mFSvWT
pTl3s4JBGG2AvpLppZWHgK2osTP9a5qPEh0NUbbsRnOvso9DFens2PZEh3iFjhbu
2dfPbi4Jn7+GlAaxTQmkwdwD3lq8oCQlHWk2nxIUh0VUtKtPmrrvN0fsodimvTFa
nneG6tduqL/NB4xdERzLCuffOI4Pglx1LRkXWczCTApWZlIEM+Z4rL9DSrcICIp8
T9EOA9vcGXwBLEOWpWSfJxpWZsJJ6hWsTz80eBdK80J1dXVWplXGojMN9UDoz6K/
KrywqSjlbi931/OKM9Y4Bmrt4MSwtHCZSUBpgdY1p0KJunxb6QVF4wE1Xq9pfCOg
UAUOD6ThUbL8h2OgnF/Z6JLLyHlyxYR8kCIdk+nq7yfWHG1BWftKUDu26yVXnHjE
CLQs1bw3QmyN7k8obmymmHv854kS9P7GobCKShFdN9kMy2jsLSuXRHXIs3gao2Zd
nFIDBa07p6YpJpSoe8tVbeltoBuIV9uGasT1QnhJre81vb8r8bMjgLyaUFH6cfVU
8rIjK2Bx78Ng1RJ2gF9/ThiqzpmKHhBJMZi5zAnu6U1rkeq0HMlNF48cOh+WB7yL
RO4MVx7iD5f6w16Dos/5Jfr6wJBEYxoIQLYi0nHI3QyPPKRimeKd8huh9HUVEuRJ
17lqhKikoz/PP2cQ2lTHC7UiufoCkfgkpFV+Fb54gLWH6jqo/JUrIfwieC40udqQ
tPAPf3l8nJe+lAZ/avePpwQoXUDEEY5jI2+LN4nd3JgiVFkfCzfwMQOmbM3DTXel
t64ia8F+TD4TtD/AcJf6rx7wnXVFZsRmPnBSfRtQVAj4skjr51tlU5Zm3aU62jIW
FoVr9/F7KvKWqqxm4BNN9Kj2JdrW+etqkxNubsD8SlKeMjOAc08lyaRECYcCJva3
ngP761P/ibV0vpiye19Mc3LavQKzwnLq33VehFXTquph3mu8AnqealIA3p5QHOfE
UxFOq+nP8Z+7WRdv4xm4bwAyYXZm2420V3BVKMeAlS+C+pOAcMJduLYi/w37o16p
EbMWjgJpG7+n1NsFUxTD6GY7Dzi22YCaeSce/cFtDqTbUHEj2HlSyOl3sHqP3PSB
DqxDqFN76/g0p+fBGVd4lfTeL5vVRYCTMT8GKsGM/WrPDNfFjmxx7+Ax8rXZE0vt
Ttx5APhUq+OvyoRDR04TlablQ+aj560yMGldPbOX2QaE1bjqrYOfhCC5YGVzjC7a
uxjYhJlAEKNntE2gNqKDDxoSTcHxyvu9nG9V57sR2B8IVqsZlPVEGgGy9DKTPFmg
IK3bjJIFwN1/p6/E84mAwfrAGAxizeF7tgRjkkXTGek9rK5OeZjG5oLJFV14YWOB
5xeoa2dj8LJJKn8Gbs8Vx7Ad9MQqSXFfuGkzWN3MxUjSJsMTK6MPanxRjGOj7w2r
t/RFS5zu8QUOMzy2cgisKYP4OleiAcjUjIcmjO4sf/PotoWcbbDgjoVSUqcUkvZk
4aoNCdALxws0PT5ARiGnlpk3sl+5rlPCR3gZCl42g09sD4J9vnoFHa8TpGNWMWb3
u14vyO4lQzLmsnFh3ki1UWr4VpzLQPabUvNdTGI2iIM24iz6rNN3uVbJNpMZHNUp
nf/QUlSbsqNacXHS+pQRuzCqG4DbDns94qTuaWc4WdOw4CmMvZRyvwjpGePCr2t1
4MtbPB0J0divVM7H0Eb7FqJVOzXE6xm6y8ojePYAEWFTD7gDA9LdUPSZf8DzhNC/
9vHmnith4pJO/xlPK1kJ0Iwsf005E9ECiDy+xWfoXuN0xjrw3+G2EdstgstEqpjy
69643P9yZL7xjzgE2v8vyK8hlmkAwyI1Tyl9X5znroTeexOM2IDcBH7yLzqarydV
9Tq2Rfy10uYiJ8PnDUntyWwLaTuRUF9kcp9AjwQttfBCpk9CDfg4ldrWgx9tYlel
3jHunGl7UTD7ybrffJONRtbH5CXl90WIeQ+bgr2TMiYfNrxdxsbqUjzeRombMi+c
txzGDc7+4B0/BK3TXuEZJtUvkeYrx7OS4ydEnpMiV+aid1RTx1Z+wFLBT67dV40e
dzhjvSZgJ/E+qfcmWYO+pHqvrFxKNoHbhnl0i7/xlYuH3gxtJjyCic7CKWqBsrW6
QX9t+uTMCRO56jKjUR3jvZGl2DyEJA3R3LcpsYa3KmT1HwaysTqovJgQj2cHXYXi
5AwxDPshH1zCA4PeEaK/MAUum67GgpJZfRTPVSGPeb/IuMVJJEf77HTbYjj5UCMI
S3jzz1k4VxSgkEzf0JPyQjNd2Wgce5FS6f3hoHCuaq53xO1mdf65beXoIEgBph7r
VRv0YisJ55V1V9T4J1YAdP2T0wpl51WLsnEYRxztOIiHjMxF6au0q5KCN/KmgUed
/64keJkR6xdD90/4l7MXSkdYLVdHxEy5TiyHC8Tl2SJbiCaB/TYgtFn+2kIOdvYe
Z81Afs8xNoYBdNJOiBQvDVwp07Y4kCuV0F2tw4p9u8qs/RzF/SdyjAwdNJI2pEYe
oPrrFIBU4BuvWUV2gYnlQJEShEufGV10lhkFi/xaRuvG9MwTErXK85yMlBjBdU4u
7t7DWaMBigOslP0r+UQq98FXh6lR4LkAWCdtwsqwCZ4+JhWOX5CYg6nJIhv6xGq3
D98DDqd0q4AewmBrT4MkGrIQKWsYJgkX3Rf6sm8JhSPwkHeFgWRlBq2RSxJVMsWw
T7USQXcvnk3smgHaIPUFlFZRcmkHYlhuZif5ceOqIs2F3x0wOSC0vAI35tLYjvrS
4uDmOAB0o5B6GBzdPHi2cshZFkC0jmsdF7LTKg2azqovqgecUB6uf0XWGfucqN+k
SKWvR062JUqhBpES7ktZDnXR5Fv2bcv7akmpAs+xZolB3eN7ta3HIox3n8lL6ZZ3
eq7atK3fuRJKs6ZPCPxA2bFJf41OKU2kLszavbx9SCE/ef6v6S3AJbJ/fMU48+uU
dm69jTBBk4piTS4KmlVtxdzb8Wvv1WuwxuNjjHrWREO9/F7sOjkPlMp6HWw0B3i+
J4tAkhJhf5fC6N5+R2EtgJOvEZjVTfDT1hX07b9J1LJNWYztMis45TyeM6sx0s7T
Dso6hEu9TR7ADADsUYcvail+Zfvq3GyaJjBTQH9nEaZSKbs0wp8H/WzXNL8KCu0+
1hgSVQxbQPWi9evp0n7QW2lY4iuiOqUcAFSqUrukbvM26G8OOxIBnHeICl6SH6R+
oFWtmPkJCp7QD90B9wp4erSU2uJ4/of40UpDl2Xw/FLU9L0gJrNXgj4L7m0r3iBT
1MjYB9zDHFgjIHMTG4xGjoGrtLib7h+NIgs71qpz49fgKJ0Gq4S2lsbyEF402QPN
kj1SJThbCJI9j5lGEvW6D2j5atbewEtU4VSKiRhf5qN+Y3fmdrB3pIsWvtWUeGEE
8FEvj4gFjlRJwHoA0Yyo/wUnRkgGLWI9F3PU4xo0BnS5FMoEqD/pomYXkQ73uJMf
G4atqR04XKRD8uHH6VHaoej0zAtdwcUHnpyqS9DHj6QmcD0e9lEUrsaCg7vJxhED
FUKwBuRSw+bfYL3/w99QbO4rrSIcJnlmFa0vgVSP9/mZqozZEUi7NTWFWcC2BO+/
FGiL12guZUh6eAj+gMTx/2rEjzbDxuHfEe839NHwNEnthSTrLudT/Lteh4a0dfaT
iiu5Ibu74fbaIfhwLWGXnFUnslWNnIHysWa/DulRXSRY3BhllqwwJBUci+hul2Bp
u/rv3LNeVxANubAQslrgyNKZBPcB2gYzPChLYbYA7l8AZdUi6MEdFKSGuBbvb45l
iFsUoUoNuowLBEWX2rgvn4qC7a3l+4UjBj+C3VhpXryNFjs56AQfCPdmV3paPUFb
2ENJuKnoRTRw+GEUWyTTnPmjfQLGZlUKalf6jgkZStjMcVrzfJuAKPIVEJETYy8o
e1uEUBbAgvF80rKcYFU8YjGROpnAJniCNLgaLsD3XS1DYzN419i01Z+eo4gTy4eO
Mm2fov44uuGlAyIEEnXpY7qglMWiOt+Gsy/ST9gdSd29GtxmOeGSUSJ5VkhBL2tY
Bq0kKcHP3Yth80sQMOTJFenYzAO1ryUJRDhrLaCDXy96e/8xydsi6/DTnMVipmJ2
r6pG9pqmC44xLXWqE9LKiuT8UrolNTpkzjZP8NV+jTSG0ZPPRJ6iOOyImn0Unt7E
psiTAbKQ9ZUUuxwIN8pgHtcHeuAOyCuy6PoYqQvga6oFGYSeA5BPdflxbfoz69+N
w9944yLl0rZdR7D+vV+fjSDRXwUHWLdkNW12TYVyMrfUr8bcoemBz4++QEp/7nCl
bpciD19vlkjsKgthbP8LYWPc3RVg3W/tIS4YnZvisLiRkZaNMc9mgF6YBe7DTuqA
Rp4OHjlVRG//HVVHBTXK4GFaRtuhOFGwdRUfpwFulqup+ke1Bqekcg37mm7NEODW
+ftfS+LLWy1FYNH1AdZaknufJtRTvc6cpKoNMP+k1R1nU1a0ijhtTNovNTt6f6RB
M1IiC34BTOJVdJNZvoM+3eyTR1lxdXqLR/JRE3G5OYyfXe8rAh3XchTlwuMvmDsM
rfIlXVI+tv+FStYeY2Us3HxYqsnzcpPwVDAJvs8Kk5AUebdMfNTfEZ1fh8wCwAaQ
cpMChmqt9wfh0UOLA39Y+/QV+wAQsUN1QqCOY5vkRyBLFq64NyTtYJrUKGoARZ7p
NDmN2WBpwQ6gMi6kMxjJ+2JAcHxNM7dDeH88y5ieasAlDhMO8l6uid4jh/GyBKZn
dPztABMMbCNNJVexX+OefM+B+0O11ifbjvToLLPy4gPIZ1h4uAp/iHGdVTMu5p6S
pAxV9k5cQfd0Ucr8p+6Q3PGP0VCAOaqmNYviIxwHdBY/DEqmj+xcgBpknuzxvs8y
GuRf0YSSGN4IZ6g/M5Uz/Ibm5BL3Pky9TeO84UZlE5StjgkmTALcWw8I/TV+ZaEE
3ssB7puFjD5GHzkNf7eyzzOp2J4dOb71j4rhd7BTDW+Gkq3BrbPQWWnleIGpVkBK
VKBa9R2MDWYZ4Cs4LF/Idz0OHXUvj372yqiCNzcxvT5kpo1xo7CBaTsCZMpTuPOQ
rHcaRQBlc+Qb3iV0541QTXuCRVEOAFzxl/S8ei8MI0HQjENR7sfAMMQTYS1xpI5/
ELxkqtNDAEV+A53RT24tMsuWi4rLWHxOhnIJna723eEUipIhjAtXCeIXqezR2MT0
8notBOKtCWI1JugbfUqL4+H+pYH8HzPOqEFp73LBYJPC04eHNiCbsfpDk1PuKGil
8HLb21hoeUahRc7cZcUD6orZLKy5Y0pSy7YaoiC7oHuCtXXxv+dcs/4FCXub4rGj
0UwcPMfAJ2W+9HQsx7ToyOdFRT+Td0CXe7OiLtVEGe9nVNVB47UbsaKLBMJRKtKd
s/NnxO0R6+VesU4IHg4pGG+Vx4hSLZC4y/KjGa+l0iBmeIxjqu1pPXDJDHPxhKzp
2sv8ODLhCTI2gimcvFtY11u7Hpuf+WTtTO2xvURYCMLEvfzZrjr1QC2NTA9VcU6h
46Td0An9MDctROoB2Le/USR++y8OWAYtKYQkglA1mIN5CqDFQ3SGUPFSLB3TRx1X
OZTUm7Y0M/OjJp7RfsaQixYSHX1pMEeaslbbLOmA2OCnxczKmpqqFkyu6Rdx71Fd
jLsbrncqTGemTEPHoY1vrgXf3LCPM+9CkRrOeea8Kpj/cn1FMkfrZcmLZd5TLOm+
0v+7K2FPNNBKfuP/kzCK0qB1iLLahfqEgUt/Wo1IhDlMIghav1R/Afs6EQSrRUXH
77BBrQwscRjB+VPvicSCjethgjkKFlVp0dV3wvUh8ksIBhSHsim8EsVNifZ4MX/K
1UJiK604C/ouVqHoYtLepRXbvvGekw9nnEmci6I5gbj9rNrQGcurAEGFs/+M+7rv
Rs4+/LQLn0JldemzbA8qZQXC2RZYS+kBPp94OMHSR9vFDpbrXoevTCIxuSlDNa8a
XHEW9KvKgs2SjeeeFt0eovylGLLC/+lJTm6g0/KLy4DhYWYbjMqdm9et3unxd06k
jHuKZuzzWmJNvm7pQP1hLgyTaAmzg4e//ja7fjQlJow9uC/A0b0cjvrpkpa0yxgO
x8xnxBG1gAT3qKdYkCnYFkoC4aEhRa6nKgry2zxK8XtR2nUohVZZdrPLn66SAQSN
fH3M4HxozwTE6DR2Tw3VIgzFuaSHyKPqIx0prPuGIJJIpjXY9/nBB6ak80MJ3kgD
yiiO6vFQ29JtI/htG74BvKuvxwXG21PBnwkGXCOaC+75cXnWW1ZFGaNk8d4YxK52
AUjZn7IWF8k6hu/KqYumkB9RArXRv1Uj2Khjn2riYsEQuSQYp7y+9bPwUUnytgz1
1Zdaqsd+18XOC+mQGL/dOvPCYCypXY1hQtPbbSlanSGwunPKbrBVB5gDFV3N7gcz
YgXrkRWYDd+Zs/kCLYjjXIjpCskpTghjtS1SADUSh1GoHLGWCJm/4VtrzoGp5dYZ
nW++tLhDFHRLTikyty4S634NH0JpAcxhTOGX7i+i1jZ4Jn63jLW0+0o/xVNyH/J9
DWJ3lv6y+HeXFwOrB8GQP08xDBuIg8f3M/tnTV2kMTJu8FrBH1W9ROfK67+OCpPf
67FjbPJJy+bqnGwOlhEIAhsQ0hTF+88zuFsv1zBtTqK4/EDPixtBlFlTa++AMno8
z2TAoRFHHzcp1Yw/S09CnY2aY9MFHkHlPDzbC7rMnCW5DU3j97mKqg4x4u0bdp7C
FAbcvDWo21SaSc4F8NwLbmPEUTyvTUoJC76Tmev/qdZhtBfra8YxQ7bMObcZ2kbc
/+wbP603Cnd5XpemttAly96tmqKVqlmLuc/OPfCdHVc9cRAk0ahOScaZ7le81/g6
Iq8z9UG3J/cQzAnzsoB0snBHOtMPkuZ/sMWg7M4z+y/q73odbGvQO60qyd3rqq+q
F4Tedgfqq1OAouk8QmTZFAwk+VePuE/LtU0RG/STHPazsRk4RDaVXOrvkBQSjLwX
co77ZLIgmjROoI8vXTh0sZ6J37R58MRSgxkZdu5H55eSgHMhJGp2SpNhh/uHai7/
Q2ZFluBVuh97RHyH4iBPMNZiJRqnN4ELhlITkB3swLiZi9P8lc7ecSreJyYKUyXH
Glh+oz8Qea39/VT00u75S7LiTszVkEMFAu26hXUHyl+bAqfY/nWyErO76cirJStB
lpyylv0jYAoj63SYyJGw0+Qi5spMQDf4eS12E+o7gnGGRlW+pzIO/3Y0rbWkN3sU
hm1WaiPcrlCWGq8uhstJthiX1mQMo9oOi+tyVxaVxS30tenRbDnbJFEWRLNLBNOp
E0GVvdKwbk73rJiIYb4uZVvqAf0HhOSnwbQvTigB2hamEV3Yh6T1WPxvhsZwLEY/
0oUTyvfWBYxHuMCSXllUROCmVDxZZW8MbRDFFO14MzUGAdiZoXihtMYJPi9xtSUo
XnjVlL31zIpxT5vcO2HD6sL0FUrUiL9MPxsp4Il3szsgLrEWbhFI1tvq/RHEkM/U
woxpupg+bjZFVE1uhK4TVPuPQjGU8yNYC9NBxepk1rZy3TCFE9iuVfyiZGUrYXBU
286nT4XsQaPiZ4bh4jVIfmb2Kbe2ADI3t2j196JJCMT1pYwClAL+49ivmPAVvvBe
tD/M9UJvKeGs8nHFQrJ5MUs44g2xdkXr2HAOIkZZGwFac7irsfnIzk0qXXl4gRit
XZDqb/lSX90sNwwej9aw9qGXL45JS26Gutv/wNlr0+Hpph0+8ijvPPqc6UkuNy1P
xYwu14iX6XzN9TUhec6FgiW3FL3+WyyiXEuajHkbiS3ZF55WA8fj5W2C/y2VyVGH
Sx1LDG8oHM5GWq6TFCfxewDkGo4lsQt4t3xGq4ofMoptH0UYEQkUSiMusfQeyQ98
opV9MN9dcfq6iF/dHDklMmfgYVUuDY8N6OIvpYU2eZVi/ohdD8Xi+csqntZ8pHS0
lGDJgwG7tvdX1Crps0J468oDD5OR7AuBh7Oz7fwFT0itKjsUTMKx9mRcQ2aq0zgQ
EVtbz8KL/k4hH5T44JJKH2EjCjTJn9lW8kt9h3QoEsoOQ8H93cKscsKOdnQxW3wq
SE88wEbroQs/d9gNfvY1Yd0DXqbZdbgax44IgpW5rcqDJyKquImQZHvqKUppEPCk
ZtulOk1lNODP8sKIrRQxeDpXicWprrWlUfpVoXaudjcxvQDbmaX6jBJiE9ufrIT1
B2VoGU9CACXhHf664Ln0+vXnJtTPtvHNy64EMaYFMzx4+sY0rSw28l/c1ISSmWKX
34XZ+FEZpdEZk3p+AzHRhj+xRcnzkTgd2u7o29SKVNBZmOaOAYQFQv2Gh1Hl7t24
lr8b2Gzk6+15u6Xf02Om0EzATARcKcNHN0K1+TlA8j/w/KqwCsudoPVVaothbQ8r
m4fNx4Hw6ym0AE3bFDBvUZ2ejpGCyIa9cG3cQbkBOnoZac+wZNuamH5mSX3R08vk
PjLX0fn5MpHW0zCs96t/s9I8+H6JEuikrCFC1NXFbv+2NRQU6hBb4q1mKVWVmsts
d2dy9jyoToCoYW3NkGA8Q9BzGcFHd42abGjN6UrYqtSq+oNeBG0Rl4y8oVVCXjSp
WwvutlUSAcNfEGZauR3EPNl9+KvCsPDl8xQygKrsgupQ3JEHmrEq+JdKk3lGy58a
4g1Io3l8/1UQ+q4QqV6hNXgp19xQkgoTdcXLF2j3fRprXEtL8/qzuTtt+Bi7PE8E
hQzM7QvgT56p+dzbLoCwIxwTAFCQHc+pvWkobAVFMc12aCuIFzBMKyoc7xFECRIP
eeuEVWOEGcq29TdIYw4l2xiiHpGslpy7j/BPP4f7mljrtOPo1lVMGE9qYl9FwYZF
ACWyt546ADrJsUb8rtXylpKqyheslILBQ0U/4LRO6SRzzCCrp1TG6+xAuECG7r4Z
sGjTgUQoKYCWTnldr8W2zcH23oAmSYHQVjh/TC7FpWfPzKPYW039tqp1xW68iCvH
vyIqzTq7GoEq6z83KjMUtsQTLmKZnNMT9OJJqjdPzZ1DcOOOopSFJIl9gU6gogun
pbG6yoi0ZnSoIqAu7PYEpuyjpMbpKVbmotXc5EuRRBeoB3j2J5sgwIEPkvEXvo4C
bfy16SnEo4UlQvsTuYkkWkkVl8+wtE3XbwKHlo43lfeHd1JNuSllj+SdKrPzjNiJ
Kp6+h3ehdQDM0ItDo1iX1hUwikL+SJcVzJYicKRGTzGtZ4DIlDmiBdfQonv5PxyG
QIv6/1NRgyXM6cyvWG+TI3h9hfNWePUzTMT2B+xBgw7AIOvcsbOPvdpv4jOaugNm
QfWOy7sDDqq6nxvw5cvF3L8OWI0XQsPeu9QW2xaNtCJVFxPd741WRuP/FlRBIoal
Ye268uSyMCPR9UL1ajcmy8IClCL5n0nQMpBbZYiO088uzpreJaf3Y2E8JBIvhDcn
eLcp6ZbvzLCHXmpFXy3euNFN/J/hCYjNDyLOYQNtzHiAR3P7hhFGRHogfgiNJyiJ
ekmdKQYMRr3fn2AjG1SR9vzap/Ec21K0y++dJcvyi3ySuHFpAA08MsRUWvBFXX+s
g+ty/gblYnxVpuxBVSc02JBJfa1EZWbIKO88qiBarba/ZkVHzk1qf/nqwgkOl2ht
+sF/Pn1U6vcYu2+94xLjbPGw3rj8WtfJ0uIi/tRdbjgD8j6M83oWp9UVBvdlWHjG
KFTnOYWSpJfj+A2Fy/lPjW3jGpJK/DOIkNqUmw3ZSvicGFuThkA6thUDhojum1kj
18kJOnETGFiBG68Hgp3rV1/BhoSV6QRj4epKwFP7Vb26daPRPiQdBgeE6Wfkdzuq
s282H8CRrhgkOyerCW1qxbZZvpIGcT7EmbB4RBd3Qqnzmoi4eIO+NJy/DOg/gSaF
8yvSoWKXp2/YKZDwST4mR1pB32S1koV82JYg4/NLf6psPEYEoNyRz86bFfiZKNJe
MWpI9qM7qjSUk+XypWDvtPiEAAVqhvntkLgpFQv5pnhZg5kjHrqifM049rcr3gZu
pkEqhAQ2e/fe9hKMjmt/aVgeBQQfpuAeeBljaGnKhrzroIwOrmti6v6St5sm2wRe
oJbSthfiVzmX31jL/Yof06rx5IAmwrH85VJyaNYn1RTXd+NOn2DOlIGEie+7ZrLl
IJD2iSdaB6roX/CL2bKX4l3Ulxf/3DHK5tk5Zvzdk8J/XBlBD+TV4UsZtJstyePd
cC+rnBve7nTWShUvvTh01voQzYR1tRut/EYBPxHjAPjhvFNpqYHyFMimPEpSI2e4
KdYQzHtwSFoyAfy0CiarcEVM79iZUqIZiqbW5NkaasB0UMmRb1Dh67i7Dgz6JQhx
xqIUPsvOafpsTfvTmc7TfP10TElmYop/XYqGyp7EKVp5ar/xG/D8pxL2rk8gsa3P
TaZIYIxWro9EHq09mRrwH7mtH40mIZG4bFJBP98qeaXA8JeUL88ytVZw7+qwoaEb
1RVRWP9jfunytnUCMrZY6Dl+kPq385EdID8abRmWdXvdb+2U6nc17EqhGwfrAoWJ
epAyhJBSkckyvtmhxoWYGECVolI64SjyiqfpsVMCi7acAYKJD8ci2poxwvKj+hlO
kuRameLvDiNTkao+pZL7fFaNRkyovrVwTVaB6mZkcQfwiK6hSLNXAPVuib45V/l5
I2VV06ChGbLCuROPxgjoDrRATWVfwBfugAyVKc5KqZoWTH2aVQD6RC6WcvGKMaVz
R+BFQBJQUWhOVbMbbQ0Fnayyry1kqWpRHxbbPV4TdOoZBKq17Tp5HORLYMOlZCtG
7PVSESvQVD/bwfrRXSQEH2hnLgD+UQjgCrsDsss5vxiF3fC9n4rkD4FTXB8rjLJ1
IMmrPjGFAiP2pM1MgF5YlmcyeI4TBT848PzPKDWdvUui+a2PcApJKTPumr4Eom1r
VscMRKtd3nUOKsKg5cJ7qiUwH46aFjnlN+AAHpQ2VOecZ1/LuCiFxExFq7FWFDd4
3tcYKGnoSxmFHXzizdMM8JzZE9/83U2byO5Sz7WFwdkwMBDNS9STu1ubEsi375vO
5PzcrRpwVt1a68tqo+LAnfklyAp2BrgLQ4zzqQZRKmhaR43vvZ9fd8/KW//jhLaI
+0Da4x35pCBct/MkAtjGnUn3vRbCkVDfGC3Jmam1OXX2j9qN5FYpFeqVDG79XEOq
psz/lYACTtoKFegO+eH2bsd9N4y9F2gN9FCq4gDL84n1Klb9/++WXt1Onxt2Zm5I
vzODaOVmGbLVEja65oHh/5SK2BgdPZhZv1YAlejp4dseHEQsoKkNYQaoGOJmVskv
AdBrY4qp6Dxsq2zYqgq1Xz7WvaM01vYjKk2GGN4mH2qyxhQIoxl/gA1TN/fevLjI
NRqFsjeRY0Fsmy4ADPeSHZdupcYvtumBsM3A830k3V+dESSpeRRgYEbfRi+fGsHU
9NZzstSWnMfSVE61vXLOG5hjEIzlPIUPxsnhIzHL0OIZJt8ud2X4Flml5Ykp2Neb
k55pD5n6LdKIf/PRGGgdvbAsB0ZzOIVkY24GEJG4UCHI2A6h/VlnsQYHal3kS7lw
g3BvF14Vci3lcCwO+8Q0VpCJwzhHEQRI43qv3H4C3ddTOyXGiDP9EMrNCzMnHiyo
WatJxXQzDBaYEfncF/ezTUBR58heKhegoP253ucexBW1sFKcHjcl0REvF5Ye2t5l
vwQjwmhM/+YRK9unH3wzvvStMWKKtdSxLoh4OSE/k577JRaR9uN7vg9r0caW7knG
4u/qllGI8VLr4p2iuRIEaqJCdaWnp+aIQX/Cdp+KBvGMWYZcbPtoL3RQfgfJTyK9
+paaMck8vOfUIVOpcvZ9vKITQovYu4WGytpINqaTycoR3y+z8kLcv2mH3K63q3v0
erLN792y3ROfxbGFXBhvkccns6U/7I/FaCG19pgMuSFSR86mY1tTUhxnn4qkrRO4
3hqbI27Eryf+4iFzxk2OifTp0wcuQ7XFnv+DAGpdFh2P91PLKZXVx94pYdR4am5S
KM9ZWRU4R4xF04XH7EvPFet5dQQhdM/FTiqlh9bzGtzr0vx4R+CMFjl1qf87DGER
dHE1M/W9xsFfqBK0+ZQjKLqtjjfjp6MC146Eco7hUsaEXTcMV9iswE69ebSoN+ns
CeDYkO39Eluc5s4wJob6gtrvWXfoWVGieQqMEHjPiQ3i7Sa8Z+/UUknDLH/VsrsX
hFVyc8+e0gX0x/IQBtQfVnhgOuFHNv3v3X/xWqsvs/wLjVG1Wv174jos4qwTksWV
qJS0koRIuLIa9rhIrm0sMQyNRNNJbyZx3/SVtsL1UaSb0JBGstuITNb2BjkbsfL0
nKBzqmN7il5SWxIQDML9fDK6DKNprEvyIC098wURnfjVI5wE+pEuSnkuilaBSFFr
LPA5bm3Xvyl+0/DFMk/kaxJU/VYcNFolDERf8xyRErhetM+c2t3EOkXwc6akmKaa
R7FNj61R4BTPoaHy/b31Mar1o8QxEAjhxLEprTkAtXh9fUzkjHu3G8TdqZQv+gjF
dxpthInmLlVtvFLJfcKpWMW4cEO+JH8TSnBr2SpOt4MfxiabzSw/+wkrHTRyK8do
+D67MJB51tA2TCIP91JpbjhQ1UW/j0VScYrUrNVBQekJfmOf1De/W8C9P5N44/PR
pR+cahiQPt/j9HGV5uFsiRR/56mUBYwrrk92A9PkNqGE+SFX4hAJ0ScwEV9/oCsk
D5PI/nOM8NdxQSpHGfNd1sU/g9XlhL08sZRI78XZQwvEKxVIrMk+TAj1ojdFP+zd
VdYVwzb2em3aRatbryvIf29bafHKmDKVYCX/PuOmHR94KVf/yIN9NfBL5R44buMh
yu0KOBFCCrdh0y17CAS5t5isaFov1xGsS/xK5M6iBzo1YqB3mNXQeVQ8Y8tM6fQP
Dq1VhnEfzvrQph3Dzk76hFBse+mYyG/e8jZ5AKvinVPJuzSYMzZSR2eIXFV4nN1j
8taV4RU2x62MV6b07fxb6hq2i8G14/EidG1h7QhxcXSWf7VKrWo5ir+y6CWu6sPA
bNYunfc1AEIaY3IcD7rHtASu/B+jg0DonImg8sFJ0FwY3F9vtfkQIEV5nQNCd74k
x8738PCe93JDTveysoYSHHo2vbSKB91TlPyUuonlbwXH05DiG5bgszILSyTbeSgv
/LOiPgfYfYsCrih1mOgtA7ANF+61HTXiAoleiyvLhT3Aqsul8AcaAaXHWRrX90c+
A0kPq9sjcoF2CX++CTuqPthN+7IiXOgjVgGFOGDB/giLukQgahAL3DfTX1X0cRLA
njsyPt7XkZ9wgcOorrTdMwIh28ARfJ/oC9EIsmFlM8qQ/J/yWiWPYooE1Csb9lWq
gubEmnjL/VW1cnlskHUI7X+M1X2FT160RLvK8AWdi1lk8wdDD9/60BC3qcrc3UXX
+Tr+R809ZZINvXBWX/BwNtyGHGPhHHCWbPGT5N6j2y/cvzaxlodkrQg0oM90NTnT
wnTSgrFbhDO23+vsC5eU7CKN/SCR6GwBdXyeE0ywD2q57P7bAvOXrq1y/i67PVyk
Wt/NcGf/Jtzfhaz/kSHdxD78SStJalfx+slcWt461dGoeBLTlg6hDdgv2/6anQYJ
vRZOkFD4fL4V3QIXIJD2KPzqIeMBMxGwKeahKl3sMkjfleTiwoW9RSwLOyJMj+I7
wutHVqN4V6VVE11limMgzVxNhn/9wm8cZFYDhO//h/hEBpNk/UK6EFcN5moz5kqB
MwPQtiwNxDQmzKDRJTOdfcoYlAjCYb6kqLmQMg4hU5jNmwaXXacJRquJ5m8+rkAU
pO+sLgeshJ9vHHRGg8tn7zv593/oszXA4HeEp+rSabyylLmxIaHboys+ZsQeJE4K
CkplvKL1+26ftALLtcMjbHRmVIn3fsQK3FwbgZ60nYUbmyTajGrptlHJJ0IQJi1T
EIvHcwZT6ttS5yZyrU8ldFK8HrIh9kDerdVUCixRvSWmDKm2RoLO/Pdqk+fh2/4N
dVrxaP2rMHN/6v8ku2/9V/F6gV9wBnSwGrrH10hEmqUacY75+0cQbSUNPg/a3qcM
Dc9bcBqVPzNB27uRBKg0+oChfWML4GOAu1ULcphbRTQQ36DKwryvFe7dynSn9vjZ
z5i5K3e3T+ZtLDea/LGnu7mQ6pU4kaRAJlw6mzmgeJw23v9zBnoXpPmqSjOJ2dxU
XFSeB7xFu6AiTkm4V1CxHdjziCZ/tlVfVUKFBHIjJ0j2eiwepshnvdCHyOw3cziP
eD8QjV5Ce+9Z9pPPf9A2R0exRm8XIokDzHhWA9L/9/esSKyElugj29coISx2WbJk
X8FigCKWYnF/AocRr3vhkAiLJ6Q/iYPlXGDKqFXchjumwWBEIfinTMgjKSQohVSd
2HmDwWIsfe6ID24VT0c5bqAwZKvVMFW15VeJ4qLDBfEpDoid9EVl4WaqNnqCfAz5
bNbx2NaGXLdWe6g1XjqoxUyihDOQ6CCmDL90fCAJE18DXY4pMQkUstsaiSEXG5W8
xvTXkzrpmYVX7nMfuaDXyXsV5PqTJjmb9Qo7IKedW/BgspV1fcXVbilVFRfr60Yq
DCxweRer4756Q6iJ8+La/xkdKw0As7YFbGiZNFQizrSwSmlVUhQDvr7h+ebRTztL
4I73kAqKnTRSc9GxTf6hry9+Q37a3Xm9Bw6A2G5ArdeqeSf8MzI8w5Pg8vnjpg+n
0jrjJMjOlwVa1x+/LN7Wlo8+VSgOEBahDiufd2OdWrkOM9tBRhMods+FeJ98bF5J
GgY2zwFlJE2SGHn5mVh89NcO6JcTjOImYBs9G+GSj5vMEO+CGzn7yCnlyoTjtnyz
vRz+TAx+uDXCXFSAeTMDaC0+5w185omJbqvmhK46XQFXpsjIa6KoylKYpw+rUPkH
HvM0cBqZaKrzfk7SbG9dJ2y82Io9G3Rturx99mYiIltUULauEAmoPZyXdWYVE7/e
f5joSFBT3nVanl1QPX1qwbYFuju4k/l5VdRdtHjLnQrrHVv5T5WANyTDKVe2BjHY
p7FCgmbNuYdZCMsbBhIumw3aPGyeLMjuOn4egPxEd+ZldFQgRQ36KqEc5DYz6n2z
lRHhIxd9h9voOUovFJWbaP4gab9zYMJWCWsZhRBnI30NfNfS0ud+/z0B4y7/HaIH
8v3OdA5Kgy3NEs9XxQ8HwuqLq3oxjIN3yuaE3bwOSkkHdf2FxTODn/NQZj/lkQcR
oEAYt8gPLsGsZ+RgktO/jhq1wsTInAj7Lp42lxDDJmaV+yjdfV7PJCPpocde4tLk
OwFktV7+XHVVXKP1LpYjCFF7r8Bcf+IRf0r9RzB3qG5iigqpwSusYYBXx++F3cPP
T/Xzj+rg6yxpNdkhjuFI5lFL0fxGp0vvL90tmCsVfqBA9wI4bUx9McAkhDUIXSzf
G7GiaKs4WsN4aq/x5Pz9aDCD7HyS+z7SrcXM79tAoRLUbDO2un6RQQaoZ9JUNftP
mzAeG+PXjEuv6nE/1yvrEWvTKDR+L9IkWhkPQnTjJOOsfjS6sp28oBPcGoyr+jpB
0NgXub2tUophqQC31oKG2J5uVMGBRivqiIWM4Ws86rCAGfhqev3Hp270CgAwJcHZ
oqQIOv9XU0Wgqj2Ju2Sr/rk91MuELPL0bMpNyWAN1Zmfin8R0ZxhC8ze8lnmDBZ/
ucGzro6PAxDixYLTLJK2DADY1JAoYhlOb/IPpZv4YXsb9Fc7krJkfBj0df4kZF/f
5Z9f/TicTFoMFxgOVJv6qshC8AZGM2MF8JW6r10jJao32o+oK0Z3JN7uyS11m+pw
/oiV4SUZtU8KMqCUaFj9WcIGj+uxHzvkj2YVV2G2kzZV09zz2ZtFuJ6DrbVrcOHG
qOoaJvDh/LAhOeu3kdx//I/G7UpecJUYV6zn0AEkCBD3Lsene9AyiHJ0deOIrhoH
8sqxY0EMOSTHiXQuG5BHnlwZzF6STRB2y3l0reTMss8Xj1U/R34ivqPE+i68k+zb
+QUYiJilZWmWnFBIbXuQ8izoOESr1CCW3uS9oq//eXgz+bZTm1oz3up5q7ICDqmu
9Jg9p2O6hXiC2mcFEEy/wMnF8xxmlMPr65Wj3CHpoHikCGaxKF1dp2R7Hsorj4WW
tljsbrzmQMJ+6OCZxCnGw2g8YoTeO4JJvBz2ubr3WC1bghFEsKT/A75S7cjUAZUH
CENFGVFgItfey5V37NuBeNoGHaPK+YF3Jn1MmvmTee4poF36vSXg7mSfFjDNhYMM
Dc1OVfw+/dLEkGR7OVAR/XmRdrYtrvZnMkIwEqFi8GS2inhpembjFDeveO+XWYNs
if7ZzZNn4QYymvuiQ8nGwy5if7XvHuSCR5379X1Diii7Vic04HmOVZlFuillo7fs
llcMNE1DGrlPV7K3WyGW41cZcRuyH0BqUNaJkfENGjbBvGY4BL+k0i5gyE5glif6
Y8LCtv9tsE+iZXmCk/Yv8gjxhSgjBCzjSOkQrAubRSUAKK8leLeH6JTX2gCrfKIj
npSw00c5O3NoZ2QdU5x8KtmGujvsF8SLQU2IphVAdxIKEouG+bfZW1CL9sc2qCuE
XdVwtMFr/jNxL7ZB9+SmImUWCc1PXccDiFJ6TJhY48juw+zn9EFqcFONAnADM6yd
iFGcBmOQR9j7mMDGeYiT5YDeInf9jyjAjBKPJGVxIv33dw/a4M7/BHFGSXlMhnSj
KAydtASouTPc7XT8qiMuiZ++rKtiLp1y0Stew1EYZW7085pFuUISGJM5QKpHSiNt
7UGn19cY7HJ7zvRA8lBukfv4TTtPUD5dKt0kLrzXthWd0xzc8y5byu2N8b7dr2Ij
KX3Y97XAEqL+4EUs865qW810cEktRBKFZ4TRyDpEm/AMLaMPl4xKRlzEZHXocExA
NtF7kKIQcuWAxGEiUwOpZb6ZI1Tj8w65d+PsQziOiTtPoV9jJHZ/ecvf3uneWyZr
IQfwP2wB2GvEuPQyLdAtmgVcWc3ai+q3k3iRb3lcgltXhmB91EPagJhuF5waBa1e
8BbE/bAZYKcNcyA6HawMn7ZXRZCeeM4wd8imYZOPuLmsBwnPRKH8d38pO5BD9olB
8aents6p6hMQshUSzp5OZ0JHt0Gp+jQs6hYw68QMnWUWVCoJxy4bBVEXvhGOBcKX
C5VGkPLtgAGXA+SxyyDPvsuYGYEPZHZgkxEVnWCpMTsXp0jJsQ042gVNv51kub1J
QDfEdAvvH2PzYZX//l1USZz4VrLl0snkLDpLvAwo+Ism2OJrwXZPq2/s2IwBujno
1NvlY3RoqkeKDVi7TNq/chuhgUe7aF1DgygCb4vH5sjcbmyc/qeEhkxhIcmUEVF2
m+Wjww88DBFpI0sUV1XSGaAqh1zbZmmcC1M4mDTMhjLJduGETOUq1QGq0YEI/m/b
AecKKTCOEBQ5AIJQe2syoYej7qW+wNmWADJZe/meT1TGLaJh8EDwjRdTR9by6X15
AlH0/3o+N/2Nr5211fat0pVwLERZz1aY8SmLlK0Ysene0HlPjJZQMfYxT0ckGYqL
xijC1Vw5WEYVhacZDltjG1OQ9pKmr/FjLGpHeaeqN/1t7BV25nYKFE82M+dlg/wj
MYsVz9adsJIeO1g/g0/zQn24LSO1n9i/Y9A3ZfcyxXI9TQkg27CC0r43FWvMfBZs
87WFlSZ2wDL4NzYnQeCi7PQvxbCSLuNwwztjoAfPrPbHtrogkWnU6AUWcRssaWYe
j374xC31Rt74OXYE3RUBDLp3MysLFGUv3lrW+6lN8T5owBvgmojmt5V3NtXUttfz
pgtW3enzWF5L64/XXsjRDtuYxoF47jocmHQnX02uM37mc8nuTTKvPb8MWxBhnX3i
VMw/72TlOG0jrVPwDTbTTYcUcSW6F4wXVrB2tLQ7g7TbYQhtiSmafWF47V+vKMQb
9w5mxew6us992uJ7iRT/N+mbFpxx5iG5yyh9uvbM6slxxlTUne10QfbHEaIj0/jV
WS99JC0ppv5/jkbIite8S95ArlRfGYUMq0LhEXLBD5Uj3IQ21zKYWoDVom0ndrc4
3waW3peOtALjfH/ts/scD1deyO0eBq4J8KzwxeP7J5xMTSVTU6YHB+jOGLV6CCod
wnPNnaSXw4KOfdfnBYM/79jF+krTjFkRvp7+X52dU2GSql6pBWJT8Sd5tKh8pf1Y
CKx/dwqmVhczLsDgLPBXU0Xee580NIIZtf0x3RJL4l2l+xf/IF7QmKjHyFZPHQPL
4qnJN2A0biMsS065Sgz/I89JKM9idqJXPMVoXTaVuBPhKd4S6BQighZ2CHHPn2vk
Z3KfDnY+XXFOwstIHm4d0Qh2i9NGRBpg/eqnyutYV7Uovo0b/ngCA66Es9saVOGX
33Q3/NRUWSOp6jx2eB6RQ1iPKFQisWfzsqDjhdeIkX3BvfkkZnv/cnDhMX2yQN5p
B2QMQ7QpDYCVthMi/9iTuOXZBdBY2yKxSE/ySXZiAhZHQlya497Y7SZPkZdr8BB9
RnciYFDeNrAu8K0d6TcsSR5tvD9UdjqDCPWhPtXr4t1ZGX+gxkwfvGqdGol7T0Ne
fYKfHqCXA+jiO+J2zU3RpIelFAgev4xPr9oUXFu2hvs6cuPek/aPlatUoHpi4sEO
tXO8vYRCGRVsnkhg5waN/HMS2+/skjgEd1g/lubUSuCKdRwOpZH6Qwkev4np4eWB
cc0gNsQSHAIEds68UYIquumXSMfkyALl0M41iLuAG4Nhu9Byta8wCT6JbqLpSu/1
qk0RO4vf+5h+IKFvU7v/IGuTuYFEJQjoXSePZVeVApdpU5NFyLLrp5sluop8dPjV
s6Bl4X+YeOc8HypayVfEJKrKODdPTmbjfsNCgkFULX78qGd0jvuR1AxeeZnyI0SM
6oqAc3eyOVWiTX7oAeycfwAhhUmACiJcg7i27K5KuI4f2BR5/G3Zgr8pj7Aakqf+
tVtbEc+cgDkf0zPEAT2uhSuKMhPJGZb/ctZiGr17Pw0SfL4drg1eZsqNxyEzqW1x
4owZS4agL8m0Md7X++n1nGG8q1gv3pxzYWFPujOxWAU/qGQrrdpYdv9yW28hm1v6
hWYnkQEt2vUJpWpFr2zpoqlGSX3xedUUXy3IW8Yu5P6SObKSGmNebeJJq+Me4KPQ
elssK+6NDI3ECzKzqQcE+DvK2QLeukHcXX6InIW+VUF+zrsc2mWrHw49uSDy1NLV
krKj+tU3iFMtpQOcxOOIf6fyqbOtb+Zik21RYDaSMhylFWwkdLbzwoCxeRgj+vfM
HvFFpfvRp5xcKqor0Nbn/4H7yg2mLIAce1VAcdpOUOyQHLlv7qYCpK7kx6U0HJGs
Ec9hOKNolvhTS7LsPGoGLSzcMXFmNKG/QR8kGIexY2MyRvBbfqLHRf1CqjWEPXdq
T9wAmJNU7oGEqcaXURSMAmMk4uiVGnLLgYzvh3PJTi09Ab5S0z6G2/iAMELz0AYU
SG4nKkDHNpwnB/0clsGSgaZfPL4J7sxa/u7aJ4R6wGoPQHj9oPd+h1kMBeWAj4xF
LqgrPUReonJ6nVtOtLEXxmExb3oDqGrb85fbXptkw1RfKKtDG74p7xg9D0MRmtPg
5unqDdcs0RcwYYp3K6vx6XU8RFsBDBrFJ5U68wr7FhIGY9FCCsBAa4iVdlp4SD+K
3t/wqrnJi7CaFxakWaljT2bKzNOQeRbUQWun1LmwfHGwgegMvDJ3qzb0Oxh0Y8Ct
yjuZOlUrnbDi4P+ugVylcj7mjyAyk4dLpos9C55/PEfAMYbQRSdJqSjh9qt+n5Sr
raBe5q/P+qDwANdLT0GTDBYDSq3jP3G/t+BJ6Pl4bpXI6jmc//LAbo3FH/uZiQt3
vjof805aYNFtQ5zizfhc9ee8lCh5DqvbXPp2x5M7q3VcGrZ6f8Un0uSxkMvuQY1c
FZsNNWhOCcpYGDSWrhNmtRiDJKVc1ZRilLwaXmI/a27R4vVf6jWScxcomkXv/ogS
/o/SjuulvRG1iHP7tOcIABCYkAgLx/XSFXhg5jLTDsFBZSPmIH9S9C2KJnV/JisD
AvVfZ1MFGx1pYw1GzpwQD1MqKiv////EQfQeO49bXQFpN5/wjJsUMvSbxp5+hMHL
YzA/N3IXBlcOfogEWr9Jg4n3mxxxfal7i4hbIeEI+7xjvX3IUyFsNRMolHqRPWBI
gQxM6lqPEJZznvhSp7ma7xOPuyDtmpt9lUCVDF3YXqNCxQWfe2NDLXEy4YkMkMFp
EKrEclNcxU0B1VWieWcO0q32/3HnpHxjT9LbK4uzCSI6XOpdPi89oxOqTAwM/d1u
30tTi5NONo3uYF1GpZVdAH3zTHXt/Dsw59hdotQjeFsbAqlkqBYJoZ4i+yNIRTcc
w5j+pj4AruDSVA4NKu7V42XUzopb/QvKdvguh7DJyYuH5gbiPQO75tLGyTw4MzMU
unghJ+V6P7Eip2q0pka/RIGHacQ95s4x+hFDuvAMGIzTv0WIo+Poa0X43Vrta0BT
IZ5HHruRnXaVsEobGxjs5AAIwQ6JjLwax6f2ywotx+t1/KAAAftiTL7tZgCUz+i0
d/MrvpRjYF6veKLkilQikpU9VW5ojnPpdNMs6ssLwqvAzJ0o8L9/AP/MY4KdSYpn
ohp6JVaqE8wHtvSxoiLCV7pSdmDBScnxgSzrsq5ovugxWu/nThH9Y5E3yw9M9VZG
HK3KPiREDqogepWI2UnDGIpV/KEN6Eb/MuK3f1WdOuIbKZnFXgMIuaPx5kSxs76y
NT2XFyQ8NvVJk29RYeB9SGr9O6A1CtFjhvvvcHCLbfXmSFDlmqiibaUd+GYl84Vu
Hd0zSzY3mUYdmZmAEPucRnfFuxmltyHA6+5MbvB8FC/Y6R/0tnayoYk2FrNQ9eRR
zpsV1lKnADH7hdBAaLUJrGRh3Wb0y8JVlQQp/ZIcoivSDi3G4RteubBY5UleWuw0
+1I0xzlvQQ8FWOboKyBUPaVeJIY+TYSU/sBDZHUW1/JK680JprrbKLm0iBmPvxxD
r/DMJb4QrbfV4Zj/zb0bGSmBi3glWSwM44J2oYmBpUPUJ77BYt3HU56fXeAzAwC3
PuSfr2oWGTus2pzzElCJGKSsgVhAobB26puYqeZrHj5FmR+ptEjzXSnez7mh1nW5
iYZOvYIS05QaWNjtqnCqFn2Frg5iuXnt+v14LwJlAkr/bjGIRcU0RpvIyPVTt/AF
Cj+Nf9lEck7yVAGeWMq2mGifrz4GGwmyhTJM1BPk1uoyel/+t9DXxjs7dt39+eVs
hnHN0OshG0OJmt7Xup7Yjaxvvk390WENGrLnq5PhgsijC+EE9Ej63eFxOPNPzQ99
dgidHPBVwwKo0UJvCHSdni2iiOw21Utihq2AcSvvROaCFZTL+Ll32pHHlUMnUyBL
KK/zmJpYnEW6dHRbCiNW1RnZZ1cxYqIVhm0UTETR1cr2DunxTjZyWAK1kr3RKyd5
iJliWPX2imFUwsQMXjzQwXymHYGb9kD4ehZXm7fs/BvkWl5J5UxV/pnIHzxAozFB
IqqZMgkmlWk3/hZDrzdaKSo/yewU7EDTS7GRsdlZZBB0DPnrjnvgy5x8JBxAJxQv
GsTtyQ0VAvA+eQydECZw43PxoAJctRgDGn/bbPytsl9TiA83nZ3pfd0DV1CyrdwP
W6MsvBnvezyBdbSsaVY3B+7RW2e1Lcwb/9UvOlLGkOOIG1dGBJTgY65kHVeOOmha
4IVqhnT/FKnCnpAxP2hLX5rdHXHHzUdePa2akJLDsxBqd2HBvEdTf1y+yyGRX1I3
CITDYUkaqf7RdYJVzNr4zbYFI6HsKw0BGVZi+GRuIpoJYFYLOAuv9JnvsgKzE3v6
QZumLGr4uXnjnKFSsJudEOTCGHhH8/6/T/q6H8NwjEShH13sl+C6b5yHfOuV3JTK
LPoEozq9Vz9T7DttanHaHDviDzQuZ0isw5g16MseXDi1+DdzCk0Iy1TXulrEJ+nZ
yAnggNIfH2+KxMnkPtiBsMvBUWQoZGwmcu9FeX8dBXwnTU4GiCqEyO8h5guQ/g5D
ltEhF+DHnEuGKzJgHRGHbyMoSLf5zcNGLrdZmpElhj7M6sG5++EbNkLcamtC1ouN
oyMUcdB4wR78JLEPqLrWzJlsxp/5Zufv2Lu1mzHTCnCNQyjQY0WqL39BuBob/yZ2
ncFxs9C+P9+uzd2jzzeA/bOjCqKLzRVwm67Wf8BphHQ7xw9gc4fZ3ex4TBJ0M1fE
3aTwCuGKuwHA+jtkmhn9R4FJY+lpN2BcdRwKgofjPko3soPstu/6GIUAhioRcY36
3LYMFEZAEV6ZgVhqF83otisCvjpkgHUbPcme16+Q+0Sj/4POFaJ+E6xi+qZvL6xS
fERQOvuQ2vCPACnbl292kI5EMtSvTvABIuod+P3MqcnI2UVLuoybdfQdFiVImsLO
Oo5STYCvX6CNXXc6idKtisNoYjV7jQ7xMLXsD9uE1at37QK8u+8ycpojUixQyzV6
nBJK9CDde/uCe8pcU7DocFGZZyvA2zk+KX8quG0nuIuagFKkiOA267Z4YiH33yST
TdjYlObIiGGodLYOeRIxOg6XL2+DR509dpk7IUb3A4kBvPPEs1mzQTcrcI458W1S
gBEB5luvttIleykAowuQKeQZHLXuzL/HevDlkDQyN/k2mgDpWKHQ+3J/Lo1fN4mp
D2qbdziyWjI8/MD8xpJUlBFYDoMrLksd/NBki27y5zCIT2acWcUcLHFr+ooUmxMk
3c8GSIbZTOEckqL40hESxbZUjV3d6a4QZMpkKNuRMenftu/5fOG1YsnHoqNpL/gF
LXb1Bx/IjIGDh4lV/nooxle7aCkC0GLECzZJk/LST2pjQcJQop5e87k49FiLn84l
A4/9slghQNgssyUWlRiM2sECty53tQcOtwLY6SCdhyYq38SO/sG9f6yUMPFGxsFx
+9O0lTExDxhlmKyatOHAYw0z4sAx2R3MXycDAb/9dfq81yYgQ/cjo3TJ28zoS63P
j3o/qpEohbDHrOQqFhwJF9CNXo27YU4Qmf0X+F/ilb34yjY25tvgNkoALZlXKBu+
SzjTnTZ/X3wR5TPIUdfxdb+BDGPthnsh7erPCzkA8/1bEP5nmcgfsQ45DjzQbeXH
d8wYymXWkSUVoHTt7BFKu+BGHwFtw12o+RxzwJGR0SAAuknKkNLiF3Jr4Tr5d02W
khdCBWM4kCRFQPMxyfqknnMX1RjokXag1FXablokjNXS4liVpNEDI7baqgrNily0
UJVj65SXfL+MyTFF8zWFBxDC9IvuaJXWnMg2BKO3QifQ2M0p8MB/yu6Ct11FnoNY
pFlXlb4NvKNYvxhyMVE/vkngwXiOxcGJajhET7/ymBRHpLwoBvOcrJmSpmH517WI
eD2dEHK8rZsGdlEeENLU43x8dXaQomCZolztJADPzsRgWC1vgmVCNguNgtv0BSQu
0Vp3cmxQoa65ZaiZeynDs9meaaWkIA4PsahTeFmkJo/bT3PzMXaBhXhm0I9wcAwy
9eJ9lQ8/dZCBOtlIYnSlGuQqHeXuyywKVvV09ytX4hgUzY3UibfrJSuflGVAwP89
Dz2dWdokR86Gv9Lvx8h3+iXozbt8kb0mskK7h8H3RfQxI2R+KgSYugm37So/+Nyb
FQAFh4jTOw0bMaW4qTNSvS5IEfic2IjBdUcf+GID6LANXX2TLsQI9FrsQ8Xo7dSF
xIsCAqx3HcyGSqRBRfG8g2PnAKknfqDqIWSUtdiWGjKuAuTavdy5oU0yvbbx3GPo
9f07Vm3uy91G5DXa4Im7M7RO+nuWOiY30YazwCMdY1rOQq6feYlhFKf5KYlw+rmj
QsOPq39XPhOvJQm2HJ5VL60dI39rX1u2vs2wuS6esbZlMRC/MgT+/k+qdbuAqhy9
09fC3JXyG918lc13lAgcg1HTGkBaVg0dxMI3nQZ08ntC8oVopjh5CG6vfUbjJEsm
KxriP/WmVbYQRnnIic2w+V0bhr+5h7jfdP9KkzF/g/NiOIQ7dpCIppoxq5/4CWJS
EAE3td6F1nv2gHGayqRTRES7zs/Wlk2cG84vKt4OLi8RH3QTNP1xachBfNcsX+yC
HEBTVW7ffQfjY1NJQa8NFJ3bZOtTSWAlo89LtX+Hemo7r4AMGbchaAmJ+3N5r9f8
i2s1Ia0mqaAPEVgswyxyBr6vprpNC1i5BFSqqd64BNf2HxIsk2IXnQ9cWTRPSm/H
lNjIQk3b3HvKfBQ4G0aQL+d9C2kDeVmvjCkzVRFQ2+VgXeX6HR8yXS9a5O23X9Fj
CDNTy1OKW/Tyd73MyhG1mLRB0vXklDvSxL74gMaNXNASDbOMMKOWNRQZouKtx5mQ
BwwcFios15v7XGF71Ht+Jt64gD/KPV48MpSBWTXR6XZF9e1rXF5hprzsqvwl1Bqu
rNdgc90RhO+261YgpL6U1l+hiWEJLgenDw6VTLlExH0xBcV4LdhPmFHLRKi8rQt4
6pFwp9fJ/MkwnkVySKtZE1H7/1RQIhgFm24LDCoYfMZQZ1DVlxVx37qN8VL3nCBL
KuMIEwwYLEkOqmaYqDKBldfO657kn6l5hp4eN3d4jV2lfWQqrE/OMjdBNUG9nFy8
NkjahogvuuZoeub+sumpCYep8embrnUuhSCqM7MuZt0oKocuNvS6bMv+rCahUDp7
YhKbBng8ESpCxm8YZAdTnokfpHvcy29Ga72L3mBz4heHc3MatcXM5I45rVnjfWoW
CmyZ2fMQkH/BIkgbsRiOyqsd/lOuYsdMuxxVcxQG9kz+N7kHxnN6Z9j4vB3iNJYs
lWwgdIIBmGsKbDnMxkcCCO2VABD6cpfADy/3TjS7B1Wi36O/TpJ3Uh5IKDOQZ0tL
HH4lvQblqS0dbH72W9O0ZOTiQ7z8o+RXdu4tB90lE39RYedscXjXyKaHpxNv98t+
6YJvr+IlKKty0Q8FqOR26sM7eEA+nzhvQtV65GGpOHIUWl8srurjBurIr7SOn18Y
6rl5k0aikFNx2OB2TQyE5NOLDeN2LL+5Qstrk6WsPBykpTIqS19ADQ/UdGyyOqGs
KDM/sUvDIgSVcwKb3RcX1Jmk2SwMQwkBiIrcNU3eE+QMhGyKtDLJs6cj/aruHgCp
O16MgxTlOK4Dtc1z63ORG52H2fwIiC14z4Z1ZC9ZVHajRYO3BIWzyuj8yll651m5
Wo6kPvUYq5VOBDBvnFI89NGZb3h7nnujczPjAe95aI5W8o7ZJp/n+IMulEA/J0TB
F0X0x6fHM+IPm/4cnmg1RPVohWU690vRinPRo5QoT7DN14db3PjVkZ1v2dD6ITi9
9E3yvDKkcAcW1icQr0jiGOTIywGGxRl3VZAvGnnq/Ykw85sI9RYRoM2LKfqvd4jL
6CTeZBkdIUOuF6cp1B2SHkUVkvbtTvz1zXD4swB3oX702aQi/N6vCiimxgCn6NKC
ATcY2NB9m0b/FzrN6FGOhiANuXmNzjKZ+nUYMnHmEvHCoaAKCQoOYVwqx2wPDw59
emvzDv1MsCCElkVGu9ui1fh5K+iVcDbUwD1Ty45c52tVtNniRZlQ+N465LisaR4s
hPuyl0JHDkB08DHQIAwzsGm2D/4nX2u7s6k/T/ZsDvz+LZRbDRD+sZm6w2ieS5Yq
GkDa20IIhHRHS03WgQymdspr8IRzBb/l12npaRJuc0Noo3ZdfRYQTuWmiX1PRZTY
4kZ0UJRJvZxoYUjip9pxq8U2MDEe4tZecX/KHsXn+XU+SdU3+gzuEKBaK9fy+l+6
HBGIzeOUNV+TmfdMlSRYwGGP8SEIKCVrRaImCl0iPx3vOSaNLjC2K92a3DZfKEY4
f4iAYn3Pefg8rDajejvsgXSpDpXvXyhxdFTW0IOK5+SFX+VPulsBu6Xd9NGjhIbp
6rLCDCN2ysIWlHl5tjG4+2WOYLhEyZPS43DIBfAtQqPRX+kgKcLnOVJtuR0BCgwQ
z/k1rGifXvBxbl9eUWB/qDWxdjtl0MdJH4sbRfRZPNc4TlvogE2VAD06xVWF0ZtO
kctXBToeosmLSYlfOJq294bIeoV7vDcUAOjv6AsWsz/Gxs+FXj2jLLndR5b77GAO
d3C2jN2birUBadgA2+ZcnVJzqKYaP8kDOIBkv1LAtDWJFtMz7Sl9D2V/HpW7YaA8
msTotWZZd3wqjhNWhaZ93isWQDtyCoqwDWnmCn9grZP7V5gkvmlrm5aYNKBdmcp+
ui4qVeXBzuud7UQA+xAhoirSEblVsBFq5D2cPB3UhJa0hE7g2uAdO/+QuQQdpzoW
rYE+W1oF+xY9bc73TEGr7wijMsoF+JO4sJRAxA/u0pwiCnQim+ocuoTu3aaXrqmr
VCwi4xGIfb7alz64e1Ri2Vj1SVTLeGSXXHJB01II06uU7HRsLNNmRVmZhXNuv4z1
lnu4DQOFcEk+25haP85GcAzKTAuFr3RqhkfzJfzbPQUIfy/pXP0qqy77+ruldP4c
ycycbKQAF4ajdvYxrIItnoilStxHX4LaLP1mUZzt++F7Yr/VvPAxQS+1GzNr7XjD
tDSgcl9k/7D5ANWe1MbSItbebfCetc0xoFXTVazWX4IAfcHfywZ/h7yFVGhZZsKy
ouKftizhD7trLnr+oIl53KAdEHX73lBRJzOyYcWLfIPDZnqv9If7HemcH15HeJfE
oE3Xl3ZiIR2aF3oeuPi5WBbEYk9joeJHsPxctrEEg47cNjLogDD0Fknom3Ux1uQ5
mEgBQEU8FcoE1NdIkaMRbIi0XUhVcgMTS6qgW5lc0zQg8WKQt/6V/kqfA/IXfw8Y
MG9/od7MruSaz+eXDmwEfzON+45I7+OH9HjftNHztwwNt6DfGZQpsya10VjMM/xY
d353asJgFIxWaWAA3Qm62YipvF4DecBovHT3PnE6lQ+SHDrsrHIltg6WjaxR+lxS
VB216oWC/D+HPpJ7wB+DLdcxhOTGk5x+3PgtR1wKL05yyLgMnLFeaON7rZ33/As6
2tUpf2ughUXg8labrzjvcLkmpLTIAZegy+agBRwAep3LciRe8WTBXQG3tzqTsTJ0
8v7pkHA7jKruuOXwxlZmRkXKWvxahCOmzx2MYZ8EdHd90U3h/+uLUQwCAAcmZAfO
HPNdislIdlf5W3ieqHeo/3SsUdBmrvOmOfm0swDQ1Xph7wLacuMEqpmRDurcV2Y+
EYMjeuO47yKfhWe85Hhgc7wEDEsOGykKaiwe/OodhzJ5d9rg82NCnm6xipN7TRmK
rsWf1x/r/WRqG4VMXcw//rIMsbkpL28cFmUY4XQZxk6i7xY/c/x38Z3r7l5B9Dpy
y+xEOALQlN7GMwJQUBqJTp4PHXYHAsmwSxmjJI+Unq4i4zS9XKhpgjdHuaUtVjVe
egKvsVHTyGKvYS2BCQQXlzGFD3MXHpHnYDYh5Ksg0jRWEWVnRGv5+UzC8llJ5yFe
/hmzgt3A0SjQzCILuXcKhrymAIlL6MFYdTxFIpFyFvnUDkJuPf3UkyMIuITE4ptY
QgmC/fpG1wiIgoZ7qgFp2bdLJdHQytOD9omIdQTFg0eWxYSgVlg7WH4v+YUVdY8r
CbSTymKIZ8+jVKgAmojuQDQ4nu41JwtAVCOGUop0kw1yIBBgXRKQ0jatDBNtEeiL
8lwct3GOpnlopSMnixcTzopdnEq+Hkg3bxjAVphUqY9yBeTZ3d5BaM6DKXLz3UoK
3ZsmkY33MELkoGEwc84y+i6Dy8O1juHxj2fSJgua0PAHub3U2ILA+xXTv8LYbkfP
eRCNHxen1Yl/+YZMe6YDlgueKMEKFnxGRt6SU9/cccbfAKdm0rYB14/x7XFmlLMU
GF2HI1Is6wFaFYA1yyRNjRH7tZe6EwgFfi+PpRU5W9F5X9BxTN+WWRdvXJjxqwPG
zO2q0WlDDQc/XJkHecSY7PiDIaI5NKdf8CxK6dYIUGaI098NKATyAV5mthzpq037
2NLsqf6fxSSK6j+PwNoCoEHnlVFXFQcx1yB2t+/lXjuM8/LsGugRvRVUJzzPfOUi
Oc8UZlI/+EpQdH/ZjRpqtHPk4ZmhFKKnNAI1flMM2KzwJH9bLi+J290o6WFsIBpC
5mP33v+W87AfxqD7hOtrvGr2srkxJ6mhYUzagL96Zs/Wg5JIFrZddveA1X/d0J+C
Fe9Pa1J6kLMmfhTaklO5VN9CsO3i8icqWn5ewHxE8IbzEHfsM+0Zfug8Hn79uGYk
DpCPoo36vnNvRl9oJVzstaAOXswt4HNQsFmwwvdscVUFKGC65NYYig0u8aePF5PD
WcVHFdg+Vm0yLQ/NQT4vmh95+yOo8MLmV2JynAcMmqM2R0J2Yrh+3hobU8fSDLrK
fqVYzIw9wh3yUJHK8Ht7ixAqnQ0q0Vtl371WCsw9DvT5Q+qz50cGXUtON69ZPxiT
0fAFsV8D6frWSFQN6vrFccRcKe3EhskwUMALE/OdG4EUmoEyRm4qzMdViwlI89fE
SPjKxsmA+nS604DXjc+qSHWu9sKizjzj+wErLUBCZYZBjUVvBqheWp89xX29l0jN
hwEFtpT3i/ApF+0murHIUIS8rjcIpEKWvkrmgaA7rqnn9HQv7nslxzYhH4501MbK
T3rNuYiIBFl3sqF7GyqFnZz3M3Y24SwLGHUVk8mtVDXRFNoV/pwXyMF3IBxkCt6k
XT4ODmxebyOeaLP8eFVR/+DtpE+q23HvOYslybRv/1vFthcB98fmEIC5/YXFpJU+
69bYkI1bzil89maToqWzosoFykM0mJCoZuwsEW5KEjBbW2R63Qh9mn3bRZrNTSdb
Jov3RRqVweJc3L3couHV0Kr22ZBIk03PuI77+xANb5uUrKoaXeHQ8aBJTMauvyOp
VRPqgEsPU9XcFgLEoQBl+Q+ugwZ7StFvGSMmIUOlIlyB8teN3/UfJ89afb1U3vIM
VENIKxH0k2HGCIHwiH6eU/Bg+eACpQg1Tswe6pzegV6A8Iev6UZ3+NO4vknsElbd
8AIQmViIVbe/Gpu2IMb6YGIVrGc6C8lDoC6aZUjIP/5V0CgfU15uh3JDcD4alBde
YPPKQFre1w3xD+xJTi7F9gQQMLkOJU8pOwNF1Fcnl4vCjI02w4yBHkbSCq2RB1IU
atA1vc+ebvckhS2RMaBYno1orSK4AO6D4LkVgI8yV7Bn/u+PKRy29dn7J1gwyicX
K15ic1EiVPtHHx6040IE7r4cSt0oISrR0ovl0HtIjQHP/k3u5irq6GhNobgeu93Z
r/nM1v8Qu238D9irotz9BG/8JiYOJTf8kX1knMBrXxmbHOx/1mjO50/3kMohYUuK
lMixjehsHfLDi4I2V8woDWaUp7ub7A4IIa1o30vUyl5JdhKOXBqPdDlF99lkBIAi
ypb40Q2fIbBx4nu9L3Q/QJ4uovjf43dW9Hb+MyB683p24JqTUyC3ZGzdCSOWlNFt
r9k50Dy4GrFveQTfa2c2gFJ38wuC48yQFspCxHQPZIEWX9JBMOqmqFYNiu9QTpeK
Wq/7YvM+i2wWeiRnJSAHadfbMOjEaV/tJ2oTfWDnFjUiNHCONZSYf8GD4Mkt0mIA
Pl+KUTUZ1LxwVReCP4GchWPU2sggRPPy3lt7m9AmCVLYo+hSJNu9XbCFmvtFi2d8
`pragma protect end_protected
