// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:33 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mvnIF9ArP5ETET5esvolz+NHPkdgIJXcBeiG/zo2uWI3BCL56wlC8++Y0kpuLC0h
T5nZHa48LXZYfjLZq/jflh+5UfQXzH1Vbj/lOLDW+empxX3TF7oZnEA+WzOgN/BA
+guldA3azspcvCX+dFjMk/g5oRSeJKL8pooFplCLF9g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 93024)
jHglqsiMUr3AQuF6lJ1gSCbNHhgZM2Z/aHX57dm0sw4d1+CtRaCjYHZ0CNGwycLH
+HwMIgntg4blUNW78DG8l/QgLqR61/r8zuj7ekoMERRAhgyaIVmVKuk8BVbAAOzE
yfbbyuSccAsL7y/mrduy4maxXz6VfKDeXxG9T+tRZ23TE7jH3ASoOcVDgwcFlvaA
l7kZWAksxNHOEmXUfR2SDRFLIqb37zJo/R4zsRWqwbFSol4iJtTeBsIGKXwkPATR
TDt5Km9Kuk3WL34BnkVesKSHn+eTGmYPrhT8RfSy4ZilfZKyultEIOZv6qIyfbjM
7P6jlmejelv69vvj1tGy43H5NCjGq9sBaxD8MbPeMDsOSt4GknMffk8pIO93vccz
m7oTCL5aAz6xvj0qCvkIqQv1Dr8FonGty5zDuez6xehE6eVAfuwPl0CcJoc2plZJ
8sRtejH2Cu18C38BNqs6s7gAlwRB11jb8z6lZFa7+Q3AfjtI/E+JXhPkac+OzERj
1VMEqtPjuBcoIVeTNk5EjVqshBUBqtggiPj65qeXz+FiqYuiNHW5vqG+LJEsE0r8
gGScbUYKIWiVhySUomO2D4O6RvZHWNwxRlv+9aZBZ+/4JCq3IFKItg1DvYgbNE8o
Mf5qFf2vAIdT8Z8O8WmzaD3CKq7D+GbGEE4qO90nJvCvp98wUZLzcdgCHXBSR6ie
vqYf/0VaIqI+NnaUkKIhdLRrvnKJTngdmKBsvf3Oenmfo5kg+AqkV+msYCScys8s
e+1RcMV9E24D4NY4k33YbLaCdcTOym411YsZG44ZWbHruyXyn8Ptj/Rk49ooWmUS
gA1Ll3ZykeW2KtEdDBNE54OdbcKBAyuZBjQhCs1/6avZSTL2OzxozLbsqyPNIxSd
yD5sc0B9zdtkMAFHk7XcfI+zU1pz8LFgYdkcFtttnKxtRutF+m1vWLQcOfTxX5Oa
8vpCEMZ8lLd7ddrQI+ozowNSKCzGZB7qVmMYkYSH9VTTtOGEYVQllbsrH7Da4q4h
JOYAzD9YJSjrIDKK0jP8/NMz1qNy5OCPnDGsbWEtLhR8GNCxTBfIu88Ie62c0e+k
mNk9mK68CCvt+3AFWNCBsmBcnQrYFGgKAvO3il3UwZIx8riR2j2CMKhS0+tTIzMB
ou/XRMN+94fVNzBECv4D1pvZanr5goMnGXEWZP6YW/lBzRMrIfYHXE1Vo2laQFsX
C2Ln19zAzSjqXNiYjrROVh9Q6ma0xUQpmbQApIk2S+vxZ7/gQA+ilfpL9ncqx/U1
SdoCmSgoLA2jUuvDLtQor3HX/4WpCBnHrF6UFzxIPnncwge1tif78zE4N8F6dHXE
BjfhEasglYlvJcKiyCwSqZev+CxKiTgpx/SOjBu/SlcfGu0q0qnnO8SaeY5uZybW
sDDZ8ucCt806hxtazemNhIAS/3CDXFY9M5HjNR39+q061XgPj2QV5G1+Bey1E6an
YasZeosv857dHTwG11OE5N8dqrU3oMHooXbB6qQ8KK7AnPv6VZERhV5dDp+A2t5f
Bgc6PGskcysbt2CsX78lUzHnc76PyhJN3tbjqV+yWmZjz6ZWRVZJZ7Hfzfqybj+Q
/yV7rsbivUUkQx7I2oWmJo2XHd6pl+1SQnKpdnIIBGNCHmKoHXKXo3wFQ41S7Z9b
CPP+V0DsGZQXFwQAfohlWQIL6aMUcFzDgOEx1Z9CXTg0SS71uatMMzn+UhPokjrw
Ib5ruVhp1dsBh7iS3YlwaMGYwmT1dh/CFkmlZIyMbpB2373zgJ9JIay4zLpOnIos
GkcaXyQO5BPgJPG8/qTh98HHNaD9M40/SsTuIAVM1Wjp+rkxorbpLIMKMlAePQSW
8hM+2xmtvrXG44+hUUFef49vYKtgaINrRZlTpp2jY+zo8vpo2sAEi5mFxj6FzWwc
pAeaVgSPklYLGL28rRhE27bkK2sGUqJL5mAvsaknOwv/Wrj5ZJP3zvezj/Jm4a9Z
eCSaeSdCLN5L3135aIOLC/RM1gpNGOFfvInTqhEZUWatLFur72RLmZCbwNEsU3Hx
fRT+m3ejrj4tSLHXzfV2oM7KXLh9syEShMb3CdszAlfHu1LfhASvM0Ei78XpEPBj
0kE5OGDopwBvaP9SxUjpmU5D0M7YBM7+tdGbx/uWZ3cgCnv9cXOrpMCxoU6aPveV
ftEPlj8XREek4DQcyZEeD0TM9QYXTdRHYFm8vl2Hx7B3LQA0KOgv+j544CWO0SMW
SMtFMCl01g65s1VzfYM2bl0Frh3KA26KdRTymhDIlWsSRZHX/ECOwUk2gk6pyqkG
2o0qHZKjo+QHsDFBAP7jcFRNd+mRnoME0CuKt75yTTi0QCLw3A9c84yNE5+/ZfWT
Lmw/cQDZMOdqd7fB89s4WbFjhNxQz7/dKiTHA+lu2vTIvUTshIio+vBD+tDRkN0P
XH2qnoducnNhQ4DNOdemYbgM0LHuBAo2KdzJ/p13afNbwu+LjVmYc2IgR/iP0pUX
YblzhebgC2ziDP87W5dmvuCgmi/WYLeb6ncUIaY9HZ1iRX0ArpbkCPVPSzFpft8Y
xz+MtkTZ+YzksL+vcAInI2Dm7Kvnkx+8o4mwQAIlUjY9I2i3hbTklVPizhQQ48Wm
tJshDSdmH85loy+R4l5z0jP9gmP9tfts6jAMcz9unfrajWj8Xy4rzigJyHHRsx5B
4FcF8pkJ5sSpRXgbjHp8JcNHsLgwk6ipYNdhhgS3P5MAPfTjxTOFkZDcY4a49Qiu
xLpVJp51r8XMLwfuwXCXK7GvldQg+kJCmEFni38Fw/OLBdcKqX69ffU682jgIY+c
fBvRsyncUQBvX49WFJ+3ht3zOqqYMVK9tuEWqiZxfqt9wQVlJ4aRPNH/l25hHMRs
2JkW1ibGuOm/IC9lEvEC3NYz/ikggIguvAxScGTooi3OqvqtL3jzBa96K3qgyMdg
10iUEpIqoSobOzcMqHKvkXZbihT4vx+72+xy40+NEeEadudg+RasLJYNpu3pt13N
adL9YudaPj1Omd5+3lh/YLn/tNqzZLxFqgmTeFKqy6UGHZhCEzFRvf1oDDn/r+69
CKOVti0ATTxPBQGJmtWB5/TnrAyft6E+UzX1xdBGdo+VWN3X1z3J0Jh8Ah/VQnQu
X2Wm3j60V5/8ribzVJQ1p+0Pwl6jrxx492kJnV9hjLIONpZBjKebUJV+lH+sJ576
EC1t57tVPSTkNPed5ZotiPWUoofnurU3v7PHYS/MkqSSkgBOJCPx8tdlIub1nVkS
TBnOazfXdw6mKLInJ+IDZKZVI5s6w4jcBOak3YlGMtBHN5I+SRTEJjUAKfw9zbx2
ot4Dp3OgVkCaenS5aWQnWH1pfoxsmB5F+6cKEeauGzUM4GjssWMsWo8f6SrS0S9x
X+Lii3OPtHY+mEoy1MEb4T7kf9uhgSPOPY4DgJg21S/BO7TNwHRHqsPXzJKG/H8z
Jzj40drDb9+C8kSXo0e2/hIiZfkd8gkpTWbtwFeoEpSDhPL1XpgIBK0pkGttOEWJ
Q4Xo2/WRhPD8Sz+uexU1gLc44Juj7kYfxN5IXYxL/QGsby2HdfPyLDB3JfobHXbc
vKdyeWr+pp3OkADxcxsHCtf0KGbdTp9tjUtqeJ0RowU0wuI0T/336Z6vSS10lWJm
2AUrBtuFd2lETgIfezHKk61Zd/0k4VhVmTwqb+MVBvpbaQ6a0RyomdooExu2Xjd4
nMhw82ZKKE2JPvWcSgRe6fzbbOE5NlUg2J4G2ZWsn7/OOqPgm4wFL4RDrlsvs3+q
ZXVOKMdPu66ax3mW09q8O3gIxGPHhb89G7WXURn7dDDVJ/tne+52npU9jOI1+XxF
TbzZRP+xJ8RyRqdEtbNTdpN7YTKwDvvldGPyxxhze8LXRce0YqlCL8ADwRt4aMLK
8srFwnOfDyhViSPGMF56IcLJQkoOv9hmNxTviYPN77cbSqMOpKqBmHpazzEJMpL5
ElWgDE870B0IfoifwlPLp86toW2xwLWn+Mqdu7FK5YpAJM7J5dLwq+gmmDVubRvr
ahuMA6EQdIMsbExoMk3Q3NEh8z9qpW3wZUCs+ntM/4S2R4L0D0thF/zD3XK7dPAk
l5SvduesDBqZYk/JIbYesQEaiY+1E2mPqsZEW/Ny/Pgv0Bpgv17jxqSBSiLbxTIl
GMTdJldgfQnCC1jJXd8m8UURkLk/uh+koBWHVN0gBkS8Q1jtagXVPOYEWVtOaL4W
KomumLJA4ewl6kp414QRALEHE4TvMjbd91cutRBYRAgqsH/qE0k2GBtKUmm5gKl+
q03pIvb4u5/aGn584y4M3EBjVQjp94qWxJpkIKKUd53rBh6U1wM4aocITn7j2Nnu
vK1WACWvTJptoqnIeodQxVRfaySpKEjtCLZhg6wcJU07TU6pHt5hHpRGqlK6G/ng
2bl2P3NcOU4zfOMPY0P0jLiSFi2xARpPY3ACTWWE7VgS2fbUvin/s/4WQjFNpnOW
d9xgVwyGwYceHEn7JWN1U8MtuCKQufdgTmSNhBNeVEM9C2qv8ME5ocZ+r7hO0L2Z
AMvZHQlt84d7djHBN5adEn3vqT759Te2wQYj282Ydb8VwrEd+ZR/HF7OnMrNJ/+X
+oXPESq8ZVYG+g2MkyTTWksNAt4lO7IRhY03MRE8nLo2+OxF23zjXKWVvx6MjOdv
z3dKOAIiVfOn+TvndtepWbDep0tHWTHGUvGq8GAhWoOgpGI33NaPWQisYvczXS9D
c9KL6BeeGWYlpNqkT38cRIIW1qA4QC/pjifHnl1Y8RYu/Lixj9X89/HIAkWROfs2
sm0ENVOakGY6YFzKWUD9jocgXyn68YzKe5n6tEkKvOBv2/AuOavJ0uN6HZ3s9VDk
Yg+UJmhMuZUJ3hRol5uuJmhfwMmgaguZPZOBRfhbfSVQJowvbca6vePijiUMrR3x
xSVD81G1A8uNtcC3EDr4p3NTOxbkSUqFCI+mz0OpyOclvdsTOV0bxLcAS2GOv8K7
I6+ViWBJiQu9z+r05jDcEVNW48wJadVmrBzfLmN9OqzfWL2LR0h8/PbEr6KL2Ox6
aWQVS38E49JA/4wUUNWifFJDuDWlimagH8DHMad7/YBguOh3FhrHpMrH8wxbJYje
C4YW1UujABQS2213NnXdk43smeSCcLyFNE1QbAW6vdpsttKjGS35cKaTlkG61Oay
gl3xTuCwL10RD3Bh9XoG6C4f+MHIhX4lNbeD60Qp6D05EGPsqovJbrvGbkOyHEqM
dmpqhFIhtdk+FDU907V0nmpkwSIY13n7ahoT0hr8bdNvYaBC85gnzR+1CC8PlF7y
R3rjCH/UWlFF/sKNwn2RNJ7swXzAiz7XJa7dKTwfetYP2sx3Vfl/hNMzJ6a3agw0
Nkqx11fDN5hPtQZP+NPGjTk6nkZpu+hOOKZW9YCBsZ602Ns8XiBWN/Cvc3B0pXHL
7xnmaMMnlqEjLmNlMqnuu80THnxFFDVabb8YmiUFtaxGTNnBs3YNYt+aCIt+pHgz
R44efW8uzxQkUsvZA5E1uP9HT1PK/I3yWXECbzj9YU9n+wVr/6DiL8OLUHl5H4N0
B4q3ykArSLQ4umfDMJnewQIqh7eDcVuIs0w7kv8bbFuFzyhDOeOyboaQkHRIinfQ
uzudCrnnKgEnBr6HoVIjivPpGYcHYn986CDiYSqj0PuYoTlGXhHrxSRzVebKpfMH
xPDuLwRon1e6VVqmygtrwwQVcW2s/PewQiLg3SIM6kPe2WIU/arqKhiDrZeAAr+3
6/+oj/8oYqD/44DXcjVEorc+EpZxZicTL3lcNlxQ5YQ4HEdyb3uASfXPNNBgHpPv
79uFJxi85q6FntP3LiWT+rzOieRTuWvLxi3F+WJL4sCrrWniiUc6xJC+Rjx7RNZl
qDW5zHUwYEXRG0vTAT7iTskWYI6gqqX2XbsSLio5Pr0hJaBN/y4F2+Kb1exQ+Jv7
ku8PTZFThOCKQuh7pvIynaPO5sMatI4oP60P4Y79MT27Q3N5IeOHf7wv8N4uHuv1
Gkh/FTObP4VX4G801jyE74zSVp5jVm7QFsAkGCpJ3Xz6w/gBbxwhxbE8dUCXq5sb
597MqsKo3mfzBpxjU31pFIEhppOJ6HeguzQ0P0kHIzRBt3AjfdhT2he+N1rrtC8k
GL9Rh5TsH+BSbu480kr5wPtNaRV4hgu7YjwOW9s1OfoArDPHjXfarPN6IIY/jR+U
E7zVc3AcxBvSyqTiFE+l2ehrym6h7UHV3DlxefjDXWT5HLl9st5bbNd2YXgLf5o+
fyHMEIvhXi+l0tTG0eeJxXYh7ApL6mMihP4EdzrhUiSJ711Sd2dxwiyvKrIqgYrQ
nmc9kZ9zZDWekM/+ovAvFExH7BwpKCEb4qGVeIo8a52OA/OGNOQj8qG3X7Q8FNpN
zvKklUvsOf+OPKL30/F0FdLmaU0qp3/NEpmH0i6QAkgR+ceaHG0G87stYL60yF+j
7DaM4AgFXOeoDZIv2/r+Gy5yvcokFwqV3Pzysagn8JVnWbg8tMWb+BOwMoo/1D4G
iwkt8E3v6F6TSS4/odNMlO2VC0HpjTPimwbdzyTXXjVffqDSypx+/RlanAdh7vbF
0eDMMoDQ21ZdxuOLR32dtb8S9bwm9jEZHmBSLc3J+pm0KoILRfSlhMLs4ad8ytNW
eMuEseqGj+0XWG/+vl3sLdCenyiBWWXSwhISdVtVvORZ2RmZVujSWdLuTg21iS4R
tafu5WSGsxMzn4O2BjfrDb8KEzi6OkVFwlGbuvcV96aAcaHoX/aQRze8/Kx5XHUM
f7ceAF+3+ZToWQteYrdCnxTnzfYMNj+WVCMaCZKbDmuNAJRHnSJ1wO5DgX3+2rkq
JkwrSNy7664p5iZz7169gwxiU6h8+PcV7RkE+luDCqTm4HqJHTbDmmhSVJOXAWh+
UI7RjgME3CzOwrtOIhOZpcdGOiD37mJFClTIG8TOFY56HHOEpoT+03evve5Rr1mr
THkOp2zJziLGAJCbfCEAbCnD9GO5N3YJc5JotFciJLElaNBUT0u5E3bTzWKXpPnB
0nuW9VTBmjK04qHZgSea5Uay5maNfHXnfX4hvt+I+IuWjmD2TRggFwC9GFDfJ7aa
gTITPjJ496IiYzRAKRvqk4ptw+qM5EnY/Hxbf+/8CPqUKp5iv7Z+w/IP3U2NZ2aC
PVtfM9UxofpDBUmm0Z2gcGSjY9k88RPiCwUv7xYmPGmu538QvXqgIGCS4XGPKtjr
AU7QSFxeOmC5krxUBIjyjToKVf0PoD5E/45C35auyxTA25bR6PVURLdrZcsKkzxf
j6JecITzY9GcNPvqb6PyAaIoc4Aj4XC3qXs+BKoiqQ3CWq6qLYMLxIOqW3GrVrKu
XrfO4lD9/zWyvPVqvvShzc4QSjO7hE5N3gc8vkxBZZ5GODk6/bYQ2CwPqIAKNfrh
m4atJgLmjv6mAb16VsgIzW40hHAKKPRkwmePx9xAbb+NYjtkEj78cwa1ynHuDHoT
AdyQFRviHZGNHuncX1gRqvW4pvO6KOeFstfdF+EpjJVbHrAXXDENnWdLXJk130Qa
oR4vrBQH831jefgrdssdZ0c/ftml9LKVkdxjsSxq3pnVDnp1I9crii2LyOkzInbc
p+C6oC6eR0a+kZNSkN6kVA/VLC+rtKqsUO7O7vE7xxgedYyYgeildklBGj7U17n5
KdyMisureQ/Oc4pQ7r18JRlfBwRPZtp1s/uEBLzrvmcPnOUa44sYju8zFcU7zMm0
HX47rIYg03RMTW92VypmHRtzMT2Rmz6XpRclu8USfXutj6rGwFIxIdyL+mJtA6+M
1ujFgZsmCcIC57eNs6GOdfY9wIgA23KfuFx1hozXQ0fM0w0zfdseV27HoIjxYVsQ
YtqqSaajCNigdtj6IwQXHLJDZ6ZqGwC4End3nH7IUAQ9OJCJ0V/QE4/2EDLqHTqR
lQH5FgZRgzIR0oY2+uhaSYfXMEqWhJpVPHFctcU3KqCh9iJD1XBFzh2mQ3xybmlJ
G97TJVTw0XHhctPgVKms2md28MIQ3xCn+XOIR4opzGTm4EkRNLN8+IDfjpr28kpC
pbYShKh5aF6H+F6U9Ewt72F7JnH0oczbrhmGBD05uMGcgvg/8SaJlGcNcBgVy+Rg
sog8sMAObFMTX5M/Yizl/cYZ4k3Pa62udoHxIWUryHr5gj+Jlllj1gROG+Oe9Yo6
FOkT4MgEnHoPI2GbC8ZmwDHnihb8yVJKSlAQElItAGav2n7RESlKaBtCkJud3mgg
cd5RzZyYdmYBUYtyO92kMtazJ+HcYTE5KDXQ8O7qCU7acQi8K6UW5vndebXR9cSv
zNekH8vyhaSnRq8yvfX15yoOUxxs6FlNdsBoqX4fOc8YjfkmYto1Tdz4im6t4hVw
2KspeqEK/mBHkE64fkxRTH0L+Co8E6r4KMt0JSZDrdujmhb4s+BwfaLocI6/SwQq
rPfexHG/w7mc7fM7c0e0vxaBbZxUs1Qcpyt5hh3bJoqsYhX98dYyptiKXGgpqvJs
JyOrgP4eIzFIWAzCWB3evlNCPjKbS8Qb1/d57iIsKoYcK+GS6ejy5U1k172a6sod
77/MgD4o+aNTLQiik9dggpof8OsEfRwKobcROy/Hj35tocTQ526CD58g5jj5H4uj
9XgjQVG+p45F1e24TfwITAvPuJDDRkG1UEpZVt8IQzbCmOGG/2zbthzUl4AM2eot
yL+mzNKAsyBPW7MopbxoPrtcctf1XJzecet15hmkkYG+0PrY81S617FsFUHw0sx0
hrL9/syIJGWJ2cbjJ0FJ3okuAk60yz52CjpH0LEmYeQUz05gSejKUpt10cIbsTxN
n2+k9am4Wu6TANcmVrg3Ft8fYwEdovVxOkNuMS9c1b1khbnAwjYAh53Y/DtoPffp
wsFY4gf1mtEtzup5O2z3gMjJgD8i6kaRO27pg9tjzacZG62fl9430Wbz1xFLd6sM
9sJ4ocn3Jfz5sutNytuHzyyUyti1+gikpoJreKfrroHKgB21AOS1kHCdcrIvqFfu
w7bjcuYBb2TL/UbTipQdx3nRFpoalLC8GOtBWtu07WWNTMPgNuxeNluxg2pHe4T7
OFBIHTu2di1OqzIRoZmjBGVgYoVr7zBJ/lE9OKiYEABUHlthP0MDd8t1PlAfbpFV
v5D8aEe7LcjZsEICV9FqQVF0R9goFb+zGz9x6E+aLP3EUuiJG6ddW6OOZAee2e31
vaEPmfjc4I8dG5Q0KcTn+ZwkauLo+fXCaoDljKuhViHFByNxJOv4cI2CUmOpJhP1
QRAAKiuiai1YYbxF2rqX+folYAtX5rvlWlcwoax1OXQ+Fi0XFnvhoa3plgTTY7s/
cCrazFcVNtKtngvWn/541Fh+d5qkSNJe7KhXwKxlU1m0fu6yxkDU5sSDY+rbtCDe
bBeT52+1/P+0L72FTGAwkUx9GozSul0Fiii7MRVLM34baaLvuGBFKEkx1H1U2d9T
8KtY4t2d4yoWie3iWfauXSXQ0nzWbr+UQkSMe25gXutnh8V92WFdt0dQYqXmBQ8Q
1qUOV0K7TmO0mCMxg/kCugdeUm90yFlIGM2aWdh+aYw1PZOOjsC5/hlNO+fUydrc
tt+KqpwOayOF7i2oiwOsMgSzYa/2FWqKKUIesF3jSAIUwArv7XcwG6TIAGOk5/V7
p/9HfBNgRyWlDzpGYPh1I1qIwKoPxyblhVV9ogarmQSaqHd8aaMZWrEkOPR0FQQ+
8lRMrf9dQzDAmt3HEK6HCyjBXVuk7cgVV+1LCHogh8T5k1yk+D0DzIwemji+PZpc
IX46yTG5CQehgqXCEm+DZ+EUkSSs+1VxMFhXlkL+1OxUJw0vxag7vk73RXS4VNrO
7rbzts6fcipuL2vbkSIFtXzafs31y4ocsIeMYrD6T9MglAjjQrISLo8Uxz2Qk11n
ftwrR4RtEAFmVt3UjM0uvm108WIVE+db7OAI0ANwH/tTSLzC6D4Blk/+dG8BlDqI
jcwetcLLe61r1R4MFlfnmetJMlFs3SGivisHj79W+ihvzYwCSCJhNu19hkD478tA
dG4g2iZt296QVHO4ldSIsKM72eVLuE2VYoWyTdy2XD1HUNNFPYxuAqbzIbeR3y0l
B1eSqUBmPB+tA30zY382v/BLvh4p3mOTqXOtJPmtkZlpb6DeRaWQjjAztaxRfdUK
zP9xN8C6jHtzdjb02nCKqsNUT1VkytvNjLC3EddVVgGo4MOr01JJa4boHLzOb4CW
VTwy763QTNn4XO+2VQkM64T+H+MxcPdba+uKZmV1ohqHDS8aDPGL8t6h4U3ixLxs
uK7yyUBLlXZJWvV/f69gSEIn/Seylev4Yv02e+9sTOV8Rg1HvRorVANBmjhetazH
u9DVmSoI4roo+LRp56kWtseRgAb+JOEbfFESEgWDoWCfeJyMWsXJ+laZh+SmcDys
VBvS2/55mbii7udjx7XJgCuyf+4yeHhRj668XwdFqLIix9ObddgY0siZosBzxnT+
qocldsUIo8ecl4Q3LOQomEjEvRbGcDqJCN+js2E/C+8l5A36FFNVn1j1GE8TFSOS
A4wlkJBYrFoDfcWgXxyGzQN1r0nKJR16mUMSCaK7q1Gwm2iqP+FxBnHIcfbwkMVw
SjsS6CuH/NLZ79JI1C1wU4oPIGdJIGEuf1yZJsrSqyMqUhRblaG11rAbvi4eQdrJ
kB1h5vuUPawWC1MZowdQUTsozLFGQvkBnNS7XuL/EXYBmnf5e+36QYPsH924Wv28
bRc1GaoJgddvpDoZJoDC0pJXGTt+ysg/CtbGf18fLMxwPO6w0KgLnQSiQueIx60v
qspwxi2w0j66gfMCbH52j2TX9nWT6LLroFg6gSDmMiJ5eY8fSt64sMV8xSKLcVUG
Urhk6VxJCfbfAdsGzqSpVLkSEOtYTD3h36nQNZdK+qSyLXHXlYwWKMZ46C7NI/F8
0erCyCTFYyi7gkJTe8deqnbCnQ0N8fiBXs+u2s8Hs1lveUq3/Qc5EZzkO8EyFqZE
FJWtLrLIDaLz0Fiy7X8TLU+clmlbdWqwJNYAQQhskuUvP+WdjjrabwHJIt9/WBIh
S3/7XApJJHZDvn+/QU718aXwkCJ+ag8ijJnUr813ZyKd0JJY298J/bV/dgNE3dqf
QRoonz0roTUThbC64zzk4GuTFcFCOZ+Gta1s/YxvbTs/3Bhg9T0vvxpDseK8vy29
xLErCoAVk/fEOPUbqFjs2i5ZkNgUzY2KPeEIyOdgwT41ShgkJWfP89SE4mQoefpu
DY6Y8+eGQEI5yFlYfJg6eDtfPnEY99y55YX5A/o6llj9J/JRveJmoPVrbovMQtrG
JVo96s4T2kiYeiIb085PPhbttWuW5YZV9qh62ej2gog3C77dY1GrTKg33jaSQQLG
EvcUXisL+kfvBDBJDuYWlDOyKULHGfEtL3r5t/+kzSpMH/HYQpAIhA1atwq5osFn
O7P25f8Um/FD8c/Nr7SlVaMLBiLwMyooZQFKwQAEvCGReaVcCsMIzv+Ies/TNADQ
DeJhdgDUcy+tndEzu2gYG2sYsM/YjdlmhHzeiDH6h80FiFSIQOBljQDGN84ox+Lr
hn37SOdnLsB0z+XIorU7iI8oqr74WNLR0988BKwRVF2Ez9/E18L91gxXeJse5KFT
9qse7aQQt7ys3lyEke2iCWnbM1vdgsbu9gILojGSX4s9ejuoyFDT/2N4HOQT9Ivb
FzVqHw9EHAXKbWMNlvyWnH2Gs9HwFkqwqqOMeTeIVXEL6KuBeWH+raVXyGZV4Rg9
cwgt4AC3rvcw+1yUoMgAsIhQpeMWpcxgcRzv4HfKKcIhkjVzluPAadVjNulvL4mb
eg+SH7YY8cTtrfaOPsjM2xHJCjVI7D2S2aLV4nCM0XYbDCYs9XpvhwrWZiA70Lzl
LngQ+EJwCYuOsARRLZbQTKfgrDS3cjPC/rtUuWoKDkSiv7bjop1p74sThJ/TKGk0
7BEVRgoE4FzU0VaWyenwNKNxHRYV4IoL43EEk3oSXqsEF6zbXiRaA2/Ip8feBmwz
Wtdb5IRlQ2w91REj8r0hxpfVTfAtXqu8Ar8jhSZdVzuw0KIaPpNhcBb6o5Guy1jM
zxbfhy/eZkJ50ZjC8z+UXCUkhtZF9h470p5MmS5d9kPGZvP7+GiLmegjs6tnc8sL
4txsddTtkpJ5D6jyUFQucGg410b17Jn0Sjut16t2ILquYCdY00wS2siQ3y6Gi98S
X4KcGOmsOBKQ6etpc6XFekVmmb7HFxD1BRlYMJrOtU71RhrYc2DTERIkAEtBWV3E
63ZQk79HjGeFvM8ch718S7AIf2EKEOJ2oa/5Iqqb6o3sRTXbtoy5A9wyBwAAdgKQ
YKzuJNfxGwfMRabLFd2gwX2cqdag1hyJiGW6Q1+nx8VSjSmnE/KSeU9KTE6nUcak
eH05zsbOLO5JtfOayZ+USrj8iZcI+zWhh1cOobXJ5hQcatfnTYZQHqr6Sh0POXnM
wW17tboH/u0EIofzs/HhHrwYHKFk4n1oA7v5q2j2TiYTHnUImi2GdNSdAcxB2E7j
Qib72wDFU1ljQwgAgJ3JCfPS9A4tIp5pGY1jEx7zQfRkNf5p8TldXGlfaOwSZP2k
5V7u7vjae09IPey4bRKZ5IGL1BG55aEQz+ltTk/YbCAL0qZtm+alegUjSBJEMRvv
l42SbIU+P41y2NDw4Lr3fFDOnqXMGzsjmEdYvKTTwtSk+g4nrCoE7zhfMCEBzX8+
40yzeHP3h7tpnD4FNoaq8nCMJzMc2bGOTwQNSeNtA1otsy5+4/KXGKlGFZ74ql8U
Pq7FPncmq2jDhJkTy61vc4MfOizrHq8uXg+yXH8HHP/PRKX8uKD+OpLRYXbFQl98
xKM8OOvylozFSSECP3IfGm4RDIAuhW+Gx61Y7FSSLQ8iOHcOouPLg6zfsiy7W2V4
88b+DP9+aT0CkMTcTLY7v4Qe3ga0M8vkX4rlKuafd8cIfKvVj+D5HAmEcimJ18yC
aTR5YzO99hPFGihhqp6rhRayBg2otB1PGUcd4jk8mAL2u+CjO6t5ikRSId2NL54G
pCzIV0vUdgLUU1SFXQMA6otXv/xYuF5ZDJguNA2CfphysjJZv5gs6zPgO5g9SwyM
7lhpM/J8Xrt5GJfFNBq7GcrytrbWrfBHoXhPaW+IyWXwaIKpOe8inddO6LA52P4H
wtkitmWBzHFaMIb1JIH+74U86fGW9ktKDujY6WOySX5KfVOUJrxzkdpKbDmoEKmg
Tsa2NNSjhfSSFo3ExaLA0CobwZy7KU0giyqB0itRzqPYc6Xc/aclMB8WZym+h4on
KEj5w9xLDruaWngVDYFaVEs7Ax8/wDeAdiuy2xV/7n/eJdLVFYrdYmmQGVNv/il5
haaHpjrVjZ7LcJfbk6Dr7HXgTOMg/NUTVtEAehe6Xpc7r7J3OS/o/kIGp+7F+2pn
zFGYJSFYcb5lRj1sa7mA+faEcC8lQ7HvWp1z87sNG6MNfzSC3eFDICdHrKVAvMF9
U1G1ibSC/Ij4BMUdOoWRqMKcBveCuxLRj0hxI5ApSDR63pGXNxYk9hmXKDJ/BX5d
uMykv9Sd1Irus+S3qk67DPwOOsZy6Qqf8BUIdP9EzLt4r8smEJd44/0LZVCU8LRN
YYLKACEP14faxEpOL3c9LZWAYm7EV0bLSIn9gxZQk2hy3l+MdBV81kj3bPgyGkNt
kIh3SI7YsYAfvFJ7dRhUoihud/8KFRDPgmoEJC8OlGTdnidAcDwpE+YuRhHuAxvd
xb478YBaIu/MbGpLEfwv4i2RYX/GYgs8OrpaDHrffPQO9nb2Aeq4pWkUV99l+oum
wuyJ6sTcPAOtwgKZQDeUiYvz1zvX2C0mn+7aFmAOIpp+eskDoGmpePV5S7vJaGDm
1913TKfYKfeO1XEy4YAr/NpiAXKTAdj0RmMvTg4KGILTpdN4qWrT7h5yO1ioXZDR
6Unmm942K294scAmaIwHu0hlHp2ooqjd4JUyyIENOloZtPLfhEvKsf9jvNEyaJFX
GoWbODFM/Qm7Kv105MdPfc3/P3o3DlRMQMr/gGGIV/3uOWMczDr8Ui/p4z5gnoWV
ZW5/4lbYdWXJYUtBIwX2pYXEicZ4caR3ZgSMyMgGFHuEvPxDw2UFs5hX4MMXe0qx
eoFQILnnM4E39Ecj10PMlie/kADLNR1eMrfVCFHGNPMxT8OpvBGRRi+oLaLUwZIt
mQJoEU4SxsCmemkSsrPIYddBn2vBqZoKUyh/2YEMUlyCNIkAZ8yfA5QSz/o6YAf9
Ghy7nypOtvM7LSqfinW3WI7k7/3Pkj7EgOXsTYWqtVcYk1kPLrzh0hKyIWAebmKL
dIcVKvo+sKxxdwXfASiSpSEz4CrayXrNm3WxjonJtGPjWMj4dW/NoHdKQmE3/m0c
pRIixTgtZ2MRxMw3xwvtWsVTVfSZG9iFPzVkAX1WuVKNhE+2MEhFjhGzp6iNFG7R
o/+Hzi7/rX7UQLMbZ42oEGJIQaBuUXxcCMDDYE3F2xI3LzE04FhYqYjAgOVWo+iH
FjLI2480cVlYj+JN2p16iHERDCREShRGM6HQH5yRMkb2oucngyU9qbY52AQMTPO+
s7XOw0zCVC2SEhihZVod1eSUih8bcWpA6l4utbCaJJ9MJLRW+PW/ra2aZAX3zdqw
QyvVR6MNuDpZ3csAaz9beu7DNNU2sO8Y9cO6/+FsVAuzpCrmm+g2xeljtj3cW/Et
S990QuvkN8WwTUhcZMMaKad5B2365RrriMtNXo7MA6Q0TSB/2Iutz+DdFgOorvFg
RyBwwrcO2t8DfXVn07tX3g03krqI4rk6ReV9p9y4eDfHB0MXsnPxz3SlYWk40oIe
kKa3O8bVXxQjlWPg20F6t/1WIty2j6Nc73v4kLU4j/I0KgOl219MuICiou8pssux
1uarCWW3YwtdsALE9QolV5DGgseKA4ZkPa61/VIAFhB84M0Y7PJufY8DFhUR66gy
Vo25Ijxg/X2klmQ9QJWaRmfxZCb6JIiP4oQq8EhMyed7UCCBWgaVKtt3f2sHVJlQ
avjJQ+YJxJ8uCIqx+cTKQpPxVsmRxjWYVopcMRFEXTwuifCc08UNyviRrn83Y9Gd
K8X4aF/M8iWA0JjJfVxv1CdifKCVbB3T3Re3mT3DMM2gNqrWrdU1Yc68r1TSO1+3
zBzI84Xzgg60WIbLe1Tk1RjUQcOVU8cHGPpDgw4oU6clr8+cLPmibGjN/FM62TA0
hiUrC7hRs0SwTek/qzouVhQ0A4HbsUf/iBRdfh4wY5uZTeSI3GmMOQVezwWAFGGK
Dqjl/r18h/5wh/e2UKJXjh7hFotUmuPWplkpshD4+DckvzuE8ZeekW4Po0ez3OLn
7WU+dCSHGNPEG4oTbnDj5E/jKjs9mll+hp8VXrao1DDf0hYHrj45V+jwXvrT54aU
tmrZ2XWDCjV22YcxPUKC5/rJDam3N4z4l2Z0i9TFhnc+MaDbhMDeUbbpMJ54GnFo
A1VXeCyMzDy6A9+K8YwJ80isEk8Mnr/pHbP26wdQniCpkDcSTgDtoP7E6SaPJYJZ
r9k9ieJlpqOKeLfSXj6L1HVTllORtaMPLjjdRWm6iJ1pDncQwzN/+6cDzd5zhLnZ
UESBAJMCpnR1KM/UaVrMAdJnDgI0Qd2Zuc/1G9cvJ3dzz86vvXPMax+9atPBYS88
j2JuvPUcMMZuwDoWa703rRt1JUhRr5xKjvLU4MkPJegbYkcsjAIEeJD1iivn8sZb
pFj4fW7P5o9WjouHcomwrro2+a611A933bDuT4volvvIqtWz0S7rOt1WOqiwJlRT
kDELl2a2x1M8WFYoIBIqursvmj/drynQ0+XocxF80NNXldEQu/yW+7xHKEqrZbA/
bMJia6s0bbA2r7KUOzHnQggLg7as+gF7mxFumxUCSjOQmS4IOCKWPPUZmFZyXBnG
q1YlsTMkaN8zSaTtYN7+Rd1tlo3Cy9HTRC1iZ7JWtc4aFzBnOn/dUyPOXVEWQ+i3
g1gw1J5M/n0wSukMe/X3LG3+ZN4ZpVh2pxb/pm/4v3xOPbGpOPjcdtYV2+a/GaEf
gPejjsL2OUMFbZdzWhEwSHMuGiI3UGXeXgqgE8eMGP+q79A1FgNcVZDpXAjgiX6l
ylASqyjd2G+cP5VNeO52xBqGVs+XYUipKZDvrjLFwa6RUWVTp+p0jsB/J89jmUik
h1PeRwZrOHDNuOQSfYnVfhuYmpS6aohhkLH7ngJwnOyL6dwi3L8tJPXCsa4BI15q
b9U8lZtyw3pqfplUzP5EORbm25SPjK9bTYV/0o/G/Ap+HnqDq29TnaRYBDI1uOU5
rdiydOVd9T6ML93yY2DtPV4zCd1K0AZbKvna3Lj41LKM2/K34WqjNxf+jOGFggmE
Jr7P18zLHdE9JBQaDqo2XjQBpVqlj0K8cHPDPmhpQGZ3l9gMc4R3ZtQWyYM0PQAq
TnqN7G2wOfnGrLILpdYlNuQ2PjrQs+xp3gCrmJqk4O/kp5MRtGlo4ongrK1VOZ+M
vzLvQuGp4MhGMcqXscdp3i7cZLerjDDPyPeYC/px8K4AOt8SIKwQ/BOMkvBl5H9d
DKnbgglHf+/ZIg6+TIOun0Tg/nG1QWK8GT4o9t5ulOwT/zyKrdpFK56YcQEtLTRe
wr7WVNrVXMUcoj5LX4fDypbwMs2U7yoAhaevmsqF0iFwmtslhTRZWwUNj/hxbwkg
+5N9ktBEP65364ZTyL+8QsFE64UICoCjKotmWAGJXJQjiKdvtoKSjq6Rc74m6zlr
W2nmJdzgiePGDxuPosbp2M3x4I/8ruyUO4hFy6oaD+JhcgeXQ6YldYmiiEBwV8GJ
j9ezUThyQDGy/D8z3lExHWmGPnqK5sR/FOB6p0z0kuBNC2iZJkxNp2vvkE5ARt+0
gdAxgWdnvvlAZek2FOXJBqN5zCKIDJxLc7dm5ChL9lCY5IWlZsm1HM6269WnMYNx
Uf2JjMAZQoBqSv91/Rjwd8lqQ5NFyhwxuhNC3Y7NJpxXK5jD2ML6v7JFLmRaFiMZ
JlQ6tocoEh7O5z4tocOylXXmBV630CjunJUywkMnPAhO4xfmLq+wMJ/dCAi00Zk+
X6SPPbW7H5L5KrDIJLQG6JI1gGzFk2QD89DsV4TLVTJ6qPO1CgeZ3sTtflCQA80m
RNeBflsSnSdYqTlNgmeoimx6FB0+SUEVjuPGzfpReco8OQXAzBsW/9GomBBzj/YW
ZQx1oY1awDa2lsq46sY24L/h7TK7AoArCTmQx9RAjnWQNgBR8+/KG8qqjcgrPan+
8oN9MC6CyPBM2dVXxy84a1dznQWcZBTjqVzKRoriD1CbMVICHZWnzbXorSkYcipM
bavbR5MYwvUa6OIZuHiBoxvNNbV1Q11BZ7uYv4Nk1OCmqVAAaQJ3pd07+rC6/drE
cwHwAWWOiq9uPdD4Exv6PL2C7kS5K85KbgScXqDOgMYPg5XTSw9LjlfU6GTIyhFx
j+xUNTS/mVGJXGoFfnusTutij/T5gch6dnbtQFd4ZeXACm6st+polVi1ntExpQO3
gBep5Ke3BCff6uL5fHpt/uKhsC+tTIbj5ae//yopv2lInbOyRBAM61I7FS7FIcXY
S8pzTILYOh2cRY/0TEGjknRWYygOQUgEoCWT/7cJRcHy4Xw42hP5bQUaauD0SAbq
/NbvZJsoK9OSnb6aEAQ4PfOVnSErpGBR/MFnZcI3kL5zDvR06IvKkcKmXPoWZWM3
EgeU/xWxHBpdgeZDFoERUNt5sXXgfVdkLKcoIybVWHsaEskDhbfY6kGI32IOg1a9
5exWuvyVIuwjENBE63vvfNEW6iTBSEnmdLqq/bsJ8zY3G/lHC9RDYVaYvHmUJL5I
ExRqJ1CgN8WOIe9fMPKZ+721C88FhJ1pDAvZMS6z2MhZqriMXnOdkGBzYHV1LO7P
TystxkhBMWyU0BlvzbroJ5oMoeZdZdF8B67myzBp3zXj5Wp4jqoNkhq0k+KD+muS
LM6hrOCUVpMhEaUCVp/jXTJgWMgv4GRDnjmP/LeZrJQiVvFfJprk6P3NkGP144iw
Im7Y1AcifsClFuZF0YbkWP3bKMDmf8grER81YymO9WQWG7r4x++G7xGOKKoLyyxX
0b3zFRqIPAfGFtL6EqBgTrEosz+DkzvQENkpvvyM/rS+NlMzJoBGqMiIO+NuAPyg
c1ghM3lE/DXUAP7acGHRGBy4lXL2NiFlsMsaZIzLTL8jAzSl8Tq8d6vf8C++8awf
p1YYXc/onOnrjvme7+om9B2IfH0cnhHERiUcHJ5irhOgXDqHEZtFatQZW7tof6tU
cO91SADp5aFe1smM3MYjlB8R403ufgvQ/3nFWNtdxklf2xTBo/sNbLd+AXazB7lS
JB6afP2THRyTL/hC2mJ/3cduxlrPQU1EDpsv4dtspQuVldEZXGhxrZQnw+OFDLym
HPpfbHUgfBfvFs2nHMB2fzuj0ynX8lNiZdEDRNORPKyUV/DPCdZWW/qwU1SFVyWU
0+7hzvJdt8hF6onvMitHvHVscd/q+e91aJCj+eAcnXXU2neWX3tdGG/XKb0/39xw
GIWRguN3VUIDQ21JkOgSMfuuBbl94/wDCAv7dmPln13oOgK6SWfiPFY/AFBntTWp
3Ji63wGAbI87noYzbXDjKkdo7JIrlvGrpI2PaCjrF7kTqP7exTG4ipJzMTEUut7i
VjUCOEPr+HM2ccIv6MbwIY9Xa5JPi5qNGy8/RCkOYQa4Ob8PKIHIfn+/AFidEfp7
nx6CXU23fhRBplmurXx5Gmyne9JnXxiIaKla7tNFT7S2KeW75J1OyjU81uXlDN6w
knfQSBvplTTSy/VV1Qru78zdyWLCp8uVL7O3sUY1V6So35WT92NTePKTIrmiaxku
RlE3CtioLxgxYDCNkfarord6lLsjv6nG3SyAdpgN7aE5ZMod4l1Bdg9bGNk3+0KK
AdEC5Li7L5hxU1Sw9QKy1BsJ/imF2ZhltdRtwWqqjwgUI9hvtsCRrtMaTc+O7c2Y
KjiF2Z1zzKaRGe3EIgVpM+LQ3mgNI0c3T2hS1uU9VEOYuA+TqRaobepTGsguoynD
IvljpGtNRwFjJMZe9Dg67EKELLYPkcdHNfa9WG/xPuh4D0XdFFydZfsL+p+Ktal0
LWEebbUgwL85Nm1TVqy/BELSK7w6Ux4zvE788KJRiR2Jig+fI3ZzGunqRXMXgP8u
dE2eia1fQ6i5Eu5SFBvUB4049zMfG0kSBiPrhXY3r0S8DnpEPDXgw3uJT1synC1h
O61Pew2mrALETafananuSeHuZgsPJVrCzi+VblA3n7QSLUcge2sNoBl/HicIFQIv
w623+hCQiiTHZMCRO546HSwSESFJgOO2A9WcCcUmbkh5fgRIBaPqxwXq1UjUB7LK
35PYbD7JKapKsIxHYnjfbHhS0qATRhgHFMFsP1xFKueEVf/eDdLBCv8jAxn/C70+
kFhebgoRJfeQypy520ALVHrm4rPD/I4Fmu7CxhjiGUbznV3skBHtW8Ut5p5kCKPo
HD2N87Tj7vuvL7mKsU6cqfiUpbvAk5ekSgPy6O8Bhydq87f3kthXh/P8PfEaO9k8
KQ7D8Edh705Fyd0IIaLRv307raQb0SIL12BTqkmnxgOCjvI+07Opru4W0aOOKxSW
1tRw1dN2hTLZaZtbadvz0CxSdWbdu8QEfNG/gTzjzJoKq+Z+3ixVYT7edpOfBZDc
iNAhNLlly46gfY68+8AT7+koRCt0cK0kfOSg35eDsDMQhHDzHLOVsMPrH0vFyhdh
GF5UUKaysrhzAdtNEvkQWHxJFCpUuJZ3lyllqY/ord4UFJWOOTpdFyKDuz9UWGRF
SQZ/pRJKqBwEdaghTm3kdl+54BX7VQCvLRxoxAWjk3KzxirOzPh05ohJJOk36bvN
i8nweGADP196qqc9C8cLeyI0It3OHpc5hrhFG1M1FgsWlbOZq1wyQam9esRJTyD5
Vs630W7nZpuYWUM1m8nr0evFNDL3uu6SSbKpjgqRwrDgmHJJOiMjllJwR99/XGiM
pA0GAXgBQuR/rd+WQqCirrMOyUtfCGCyCRBgBCvWJH8QTIKSXfQZO+0EgXOZs74r
BV2q0Ej9v+iefoVSnDahC5GFLYBh45yLUcu1UAJmvQ85dgEZrI+KdERW0aet2adh
/IpQi/6uneW3w+6GmtpLyXOkwGiflXtK1rL316Bch9LoCpUsjPr+g7Jv2zdhu5mP
yMyDz658eClzxF4sJrB6ds3tRbxG/IOpdAG2+DVIOlpbkm5ndn9fL/HCHaGuH9fr
PUiS2S+v1atZBgN1j64+6flM77mmiBzEGthoRcbAHWr6ETDv7YHdHwAd/mZcNXun
VH+UzUr1IysNCqTTWzhh12Wyw/f/+D4NMNbFUymY/e+b7ppJ+mS9GlPEMLGqzPG0
jcW0fJMA7jFGLTjnllPh5jYLaAEk3JVlM921MMRxYBs7CzAsv+PNSgZPiHOCXz3B
xiHtgaG8UBrbRQdh6D/NgY4fNkCGKtAnYjTH5O1q+UiO/LZO5Fte0UPiO4a84lzQ
aOXhyyZjQgcYjjSGVjpOIgy5xfc3eackVJ1FLtxMOAAnJrkGCgWLZxViZKJlSAIM
SErKINeMHDREHfU3bG8EF4znaQHU7saDMHk1IZnF6JeAZFM6/1VxOOGGcuTcKvqm
oVSkSqeEErCjvMHAVJiv9je88XMzWm33cs18F7fodCQvcIbQjwv5s456xRU9zUTk
MSDEUyzXoDqebx4Hz/XlbQT0FyAmT/b+QQ4v5RBmMJj9RkHHZZ+9y9nH81Kiu4SG
ZoQ5zK8y45RYjceQDaP/1kV7+fxYbdZlmnpKRifsdxcbjifvys1kMRjIFE457+kL
zfJJ7XV8zYPpSbMNxeArt7wtITEBCwXVQFy40CHwAGzZILL1SEhAQII+dm5DLLrx
Vm6w+PHMx+/TocyX6MrsiF/yt6LFlVOpETKiIJu/jNfVo1iWGNuGeVWUil6KowpW
slRC2h21yF71A65y2+t5L717HLTKNLRnUoi8ytcCnkFHiYFyJBuCahmOociqSbvt
iPqHn4bv7wwxn8vKUZl3lQrBxFheOrlby3vTWjhb9cHD8adYYVqhmDMB/V+1KvpT
HD/gVEejDAf4cahAqeFTmNaVP7a4GKaRWNBGQdkIyXXIm/tmiFRDNncw2gaV8oAF
r/ldsx9JG891VNwSZY9cmKtQVgJZjWNPT4BBhCpwilSPsWzdXMIiJQERRIzj++7c
kD6nYXTqsGWqXz6uHVVyADWMevd8j94NHVTp6RkqRp+zlpgqBjxiTAt9ZKbunrpw
KZJGylTu8mvttUXbtHDjw/HSNGQlqNHqNE/vhyBhVA9mAjkEFl1iYvSFcV/wks8m
8Ls7+v8ZQSsocymQ9YhbLUWZrUXDqSUe191AkiBxC81K6LZZjXIyaILNOZArcHQX
aYDbxHABG3/MZz3/2U0p4s5LuOijvp+BiHWMEbdW4ZL3/5sVuBHpWPVTOPX2v5cd
DLjE+jdxyNIYW6j8zaTmUprsc5OXsrEo9i+ANF74rRmnTd3/jiF+TpMq3w6iCUB+
y4W3RurZuqOkiVu7NjmnVAiNWzbY1d+72QVe78aR2yLgJJPUIrfhcnNKjnApiCK3
4bwlgHo8VS9JX0+7wMO4sjUw+RKgBSGfMIIFCakjc5S0waII/v/0dMjhuWhftiFC
xzu4GAjV+l6Y7STfm94v3UH+3M2K4sstPQhwU5l/PlFOaqlUWbINpj5Dmtojsu2y
G564bzIuH4cjfmAnNEmgYpQEtYyVpOyQW+Ao4teGwnHlOArnn+5iqK/4aeAX27CT
YCfeGGPqkhqDcXiCeCwskFmkpUo8qIFjpGjypj9W6edSeWjKdH6kSqKsgg2ZFTJV
b5Z0OTf6vbWnxyBq0H+S/7ligh0+i0/G7ANPtmnKqRTKUQ9hdhLrrpnU8XgkKWn/
RegniiTiH+wx4K4giLTVzdVwwpeUzf0BQvYWCIYEsFpKkQduEuswo6jMoqeAgBBU
J6pFrj2InThHLaoHlAKj9GFqOzler8mjTlzsZ3WlLsWyquW1qUcLr49SMhTMVOYL
eVlPHlSgNMcEQpH96QyrqQBuzBx48SGQHfyzLK/7wo5P9xsO4KBYK1t13dyGlPh/
iLZ230fgg8MkTc6SG6TwtgPfBc/s7kMH5dy7M7RKvc+hko8ivBZzDeUsKh9oza/v
7wLmUlWS4AVDHnuywN8WzuyiCtWq5d6NHMgMcsqyIiIkdCTWFyCxaVIzaTe3SplJ
OasJuwoKiQ4zdoKqBiNZHfki9Tx+xlJ1Vs5qrYIKiBILeOAN0+ovYyLZ/u2ZKsUc
sIv7E7fv7Bm3sYTiW6q3HAZmyj4E1I8rIwDjJtaonvWks8ve4AwQDmT/OrBESIpi
tW8mxtuGxn9VhIW3kPDT2AdQlPrqboqe4ew+jCZ2g6zjRzhg5DbNsZdViW/dS9tg
2b0N1QL/84jUMkfESYWUWt823dr1XT1coZDZ/P8QpX/RUO6+OBvoHSTLgUzH6xW/
qaG2+ZSNCdqUChF1o5SGwdzGBeDyNS61ZaWXbwrrNcDLp5ETPTuayBLwaHPNh0Wf
I2cKO2BctkZk/abmc2MUIAa4qKFObyYyOTfZ12T8Qt9+OvY9fxFq7bOGFp+T0g4T
qfFXZeqIqeeH04mz6bdo0fABZG8EUYx02PQVV1dXl2xYDcnNHWtQS+Nx3xPrAKAg
MpHGTztKIVamRA24hWNPi+sovm4KNOUasOJ7dbdzsTSaIJMjE2f1lRSk3mznvTqR
pfHqlfHQxaM/JIkqph6jS7jTt9ewFnJKjJqhGbnR5DBOQYURP4Y263qWKj/WCjUR
GX6/Tfqlua8Z+pqKP7bPssXpKjQOkp+WgFOzu1ag2baEKuduCYnFsjxV5sdWyIP+
80eM5jNq3P+d5hAu5Jg18A698hmO2Oa++zIGkebXsumnizag/M8IsF3DPMgmHrWC
VPwXcvBNrRcB1qGCJkB8DJ4OLkxdOhMOM0lO6Xjh0M8Pp12eHDCeTzlT44sRXCvt
w+eNj9XIm0xKbVY9f5MjABgLJ6dxy6PekVe5H6RqRSYVPHQ9GstrzKUngrU94dOv
VLw2Fv+wiL0uqz7k5FYwZKH6/zvUW0wkJS2D6bWNKz2KdLOk97XoTFcmvNS9nzkk
78wI46j3d7ppWPx816EfOhQYVCIXZTHOXXCLqksWNpE/u4bUYC7zlBbWnzBq6y4t
M95LxYX+uHRmqpeoHHTV0+CmliCOE7LXS8KCdg2ZpF1V/OaowgqtUfahNGmWQjI4
jzaVti7k/CU7E7wyah04o6YcM4Z1DNCpx8pjAsCBA9cO756258Z8A5dFQ+xERI8S
SpSGNS9arrRijnziKW6ko1rtPQq9vc8WxcAhf5gnAxIrhQsXR8EVlQTJnaZ3VkWS
BIFy4MVoy11Gl/oJqwvpRuBxQCl73fTEBAnSMrcElhQXwdyBQdsjgH5bEagj5okC
Vnp5AqQiiSud77CXGM+f4blzXFddD+r+MgOnQTru/DgUIRzdnt83X9lYL67oOQBm
YNP9DplM+4Qn4+NCcg4jXPumdzpGRdO8fpZc5jzoAMpayaWLKibtKj1tk7IhIlEJ
bVL46ABPUV7UCd+oK4KezW4l4tOBHIVrZtCTd8vb7QLK6bdTT7J/UCskOOwQdtM7
NNNERHaam3BPtvhAXKySZh/xkQTwqnPpfXNpDGfx+O1aRqA6HozKDtGIs7YKdrQO
tV4qI+dCuAsine/Ftf+ce4uqYxm+5EbBmawcd7KZkwWxTmY6BENqlUwqwuCd6KIV
dxI17V5el/pinuiMjDfif3gNhSAdHPrCiScw8E7paSO05YhwTWhMHVinNK7LLBKu
MSrlP3GXpAzDLV2vGl20moT//HafFFsCDNOPclvUqsyVZkDumvapiah/02u4ebYM
SHJDnhaVowc3g5El3Rmz3tEHYQ0+HQGJzVngBn32l4c9FXJ74syfoq9plepeh5KF
n15nloGV/h/0KtEwsh11qMiaV96u5GtMzrgbiieobz7a7zGsu0huY5N7VmFhTw3H
JM14nbxvfd/CRW1RdXp2IxnWDHjNj8RYHcE/YzoFpIGpKaRiqqlXaltdLZTOw0b/
z87Q2LDp6verbv7w3MfQntOwn5krE6CL5fBAPm3xyhjp1/wKfMC6uwPePoARm9RA
ipB9JM43hv8Ac+SFAYCI1luGy+ZbY7oVj5nNkqsVNB97VKDUVdAlwzALKa8v/pbE
GHe5MQLWgCikz1PP5KjKHHaLR//8yFk2/enDT6BpnCdZILZPMdzLvW7HaKWBQdWh
I5DaB6YVZpmJiK5fq/wE84yTzJ9kCp9tpuLsFJvIh344sFjxQCaNPrIX5wRcFanv
u/E6B9zSU5V3fuTmC4g0H4U+GL0qZDlQo5kr+cKKXgZi7nn2gYzNwSWvt/PSE68B
WrIPia8LaD+HtliaCeuSNHpu1p6E6T8391MNDrtg0Wk0mk5AiUXl07nSyxICXS9l
+znvhxIPOBp9sILdpyZ+y39DBL0vkJhbIQgK2emv5KDKV1fUkpYIGWyZo8LlPJU/
ePwEP9qCKp0tSuh3Ngdpne7BfYka+HgENV6eDOvi7SSH/6dMYy92wYojft23ZpBo
8js4bGpPxtMOBGKL67UBddGQo3QByCIhn6Ap7bosXnK2OJ9i+3Bo3sKtGGEKEH8P
PjVPF5btHImn1p9ONVe4nn5cAPDA9cxHThVWxU2nRDaohjNI2oG0WxpWwcPqGmD0
oNc+lOqKGzKxdDA2+nbUJTrG9kjYcNU3xG18EV39wXQSOxjmG1302SWBHMw04hsu
nJF6ibo7T51L4u0MXK/4i+OTS4oXnrxF9HQHTw4keGWpuHyNCohzz72kAnsowUbE
/tJvhJ5nnxrjOsNvEEAu1fnIwVf9haIsPOx1jIoJ77jhJ5VgHKeVua4+bpTaFNWo
JWn7Zsq7TC5EO3cMeko9poQvseJIF+3EHU+O2VjKHWAKrSJPcDvjYA7pd9/dyvxm
uEtomtn48klFL8Kq9uUTGAkynVl7M9h7M0UwSKSq5Lx8W6hB52n9m2eouv2OZAdw
YPO6r5EAJnfF9ezVzw+WWUEBLHw+uJtQ2osLBzojgjn2iV4urttf/JPL+0gflsVj
k0uj9qaa21Gz7lIOl1otzIjxOOpP/0TJK/91/Tb/BLyXSIgEnZY0F+9IeMk3ARDc
KN+DOv6LbRGWxK4q0dmzEuopdUsJZuTfSAlt/kGwsL286PF0pk1r62/r60d4VW9g
TLNUU0z/MQ/YdV0Q5NwERUT4chsU1kA5GDTNJuuuu6y5ZPtw5poFxSKzwG10etii
5W9BWeU4va5cCqVAGmH9nc7W/JS46ySZuZYZCgpn2C7fufpsJZ2hEsBmsXknqQjf
RggwgefHebON3jqRI5K1rQdfCX7XO4M9AN9yp3xcpAUfpHDb3eaN6p2jT0NbTZRI
9oPKRx+HJF88NZYTjUhCTpSKPQ7fi80e4PNaPuRgYulvCeRsboAqr2YgB2v9ZgWG
u1Zyol2g+uRmWd2xig4WBtLDjzLSdwc7bJpPsyWWzgEzLAalp8l6rThziSoOe3f+
gO/HMym7yt1ucOgO6F/f6vY9lWRoBf7ego93ygMo4JrOYLuyc9xOoAF+2RaDy8Dh
d5zA2K3KdUYUJ/zGSyGK/6DJVIfc42Nn0z0V0m15bU1oSh7bkWYzjrpYplER7BCI
SqZynh0tF5izXqDln3HAT3SZBs23uKaLnD9nzWpXwg4pIXemeZCyNtaZ4m24UKMM
VyORnrMPZW7IhfTeW6ucykYTOfuSOWkCtFStTOQFbpA5c+5KOTTKrA3zrRtxMppz
iya2sQElxDBR/OO4qlFUAp3Ap6R0ilGa+Wc0fmIe7iIxDqwc0dY5EaZW2Q/RCps3
ki56PhVqtghdHRSORPwohSE/5J7klHni2zFEoyMIM9RacFFDsJmSNOqgP5IjbwhD
EvAoOYct3ZPt/6+/SIIHVKnN2ybcSZ5Z/yIXDSEQBH5uGgm3Xzh4AFdhZC7WEQh/
SnWOD5cHqhx/HKvOSPwKSev2XAJequMQP31C1zYNf8PobocfSdDgDd4ODg5EVOTL
3AFrBO7PQPw/fVdlrnei4p9SIo81l5+cMK/uKzpkHpS9gdClrmE0HyFLG8yyek3I
4eGA7oSVgr1VnJccENrsZ0TIajiOCjJt+ZD3hKTy4eZ2i9p00qXokG9g+9FwXR3g
hVA+MJYHZx8wX/NxNQUrX0pljnpc1zSQv3Omhn4QBi+FEXvibkkAaRGc3mj7/bXg
NCTHMHp0qQ7xQOElW0ze1/i83z5bjwGvf1YNjMLAjbv/e4CZfrY+pKeK+WFHkArL
fOjMSRZbnFrFg+chnyTJiBGQxrEcH0K1jvklGkA6Wk0jTpQTiLta0SkTdtU1DNZz
xHDRVZqKtu8XWksnya3HPEnPCCpZ22FCQG8BMpjt/PVo9+Hl0BNNUuyJ3yjMvd7/
20PuABS8j+J23Q+W+ydL8FF/1D4mNbP2ZcJ/tg2ncYocivWMmpBMJGgka/qaC141
5OZDcmCnzBQ7dUFA6JE7845KQ2Glu8GjMG6dklux+VeIt0oejxUzSNiXbpbhpLKJ
1r06MPdf3PTgE+ElRZb0oyroOBIrvFLdmmBHOWIXyihehY5Zh0Fg92Z+vnmfcs+J
rm0G2pbKrFxOWg/yno9gU0Ebw2FYiDDvBNQagDWy157UH8AMrCTPNIPNi39JT/Fb
g8UoEIUDrSRVjl+X3iA9CZKW3o6Ewx3enZgLUa4WuxRJ2vrEltfxH2Az7rz914rw
iKYAp7lo/GYIcpX6X5zBpPLG42H/6YCjwpz8AIUFZR+tDZBbcjTZXClbklULv8Bq
lYz+9HtKb/PNYrBUF8+RJHIJS9DvjHym15JDFxPBiAqNWPBIbiKCa9xg0ufTr6/s
bDlNb6Cw849Xa0OThd5EaxbO4IKBxdC6guZHjBdSGuLZmRCe4mQNPAQXEX5XAzxS
qniY6CYeP2+h/RmyGb1us6hwRWxuDF6UmRiHNEhVmJkFqwxMwBpItheU52Ss8Mw9
xdKRRyHLuQotKYQ8EJHnRuUQlqn25rBpWzvN/axdOqjK2XzNW/SWJ0n/rbZATwnn
rz7nupSdfGaIEpTQbv9PO1sKT7aPQAcMNzL1ZjPqsXHWskdQOmk4LWNVRs1yuVzA
wwimxwFtkWVpaJeHNRVU/Z9ZXfrr/0JOe5rh3zESW0fBrrVRlDVaTYgaboCiOxaD
LX1bScthlzaFg1BP04SOead8HcWzerO9ialfESxLBWiuSnUKOlasyEGce88Hn287
ROlqM25paB3gOCZXvnujLNS3RmRaFMWB0ntnBmyE4ScP4RlwBuF+xAZoYT9NDtSr
HbT80qED9seYOhZ2wpoTL53qnmykxaXosoq1NU7gZ9ZpeCkTpuRBNvkcmP+YwPXc
ZZHt91lb5Atu6RP22FajZ4O6HW28nzuUjkV0QG7QmvuxgvTk45rg0Bn1/h5ObaXJ
FdeP71Sr6oOzFkQ5ovhX/wzKP6qqqCU+B2EsJJ/P22Eh4zEoqputVNh4mmXjPjUI
1wHoS12R5SRrV8GKPaPcuxJvl8DZsS17twJrGi4SsgptWMhLNlHlLjnRW3O2EM+r
A+OyQDKGbceWjRik55rpNr7PRrXZ4HGxmTOIoO4htNc+WLwyVA+7l0Lgxpcu70P9
wCjvE1hnn5toH9ikt+miKD4Qewr7uQ1qX0Clit8JkwcJyfEnmsOmRzBkcgSuyhkr
f0Bk0r+4ASuttu9jV+DIF3aTe9qtC/AHm52cvzxJez9Z2O3kxCcb22U5cJQDG9da
1xmaJ54uAcVqwWsCgEGBunbd0pvv1hql8WHy4TT8keVAjyxoqNX5UX3qoJPRo1WJ
VN6H0UiMJvy+jg2aFvFcYELdDojrcbXh/7FLXTOyM0JT6jsuoK7sbl1SHGWGdJpH
Ap3bkIzY+vrZXKfXrA4sdiFZlnSKhrJe1RLjkGbWxte9g5/h1Oe480pKLWWcNV4D
mEHE15uOGql60IYhfWuQMSGf8Bi8bnsALnop7w4F2FRwe6ppAt2ZCT7HMuWkAYYq
xOIX8YyIvmn8lPu0ZMBTiDkySP9mvEqGcC4cZ9yKeRmU6gbxJLEgXNmNf9lFQNsQ
rv0+KqTAefEroFHpvqJmGbUrt6T4Mwm29o66bfJYuDhWfossdr595PdN4woWKZVq
eXF4Oavq7OsAjoePXWeK7fMSKUvehymY71Mj8TduwSaFm6F6ul6IqbRAUbsp7wB4
vZS1k/03mPHABILjGc4go+Jsz12tJ9NlTMiec3ePv61bHyr80kQHiEjrhEJ1IDcy
rxPwuwJqoTMFnpIKI1rep35ZSdyJ1XV6t0EDZ3WWlVN5m9vOK6/bRbX6zkHnfjn5
eKcCttZ4lXy/CxkxltVweh45F0+muSwoaTWMTiFGeNgXPML6qArzHRHrBj9cKdMa
+VvdRnEecDmWe0yMpgj7RhFblctjiMmorpRtM2EanaiiPUaGSmdgJ7yXuYlAAZfE
eaQpULsiBqQzyh+Jn70IhrfZH5pUAAG3E39Oc9y3gb4kcRy693bW7F3m7E9JGWZv
P4KtmJAbiuMu23dRZHZrUshdbAutXOs3Cb+wnlwPzWyDVzhjz+vDBWlhJQZXE0SM
6gPbyEHnb3dX+wAClk7+sFJlDJBda4GmergYpqduOXtdT2kKsTYIWSAXEHBbYVAq
+h7wzcBfkmnt06nL6XEy+DpzcLrOIISkKOhNQ4fnOv+IMt57XEKmDFs4kpxIm39z
Bks3XxYVUTqIeedV79Xzk67bHO6Z8BlsHlb+uZPpZP0yPjgHYg1SuD/UkNf1ls5N
gST+XFAhr+hQCI4da8Z7MY8CUIpNrTGXPALe/gm4ViUBIQsURBp2HIWmzBarpQrR
k+KN5wz86kaxY37pH1vtG6+5WYXmbDeYb807/BSHdcV8oWwHplY+kWCarMn8QiH9
2rp5wV0Q+GQp7O8mVJ5mbsaCgG/sxCQIF46aob31vAfjM3QuARF28wUFROljl4dN
asz0bxsAjuikvvvkwcTcIJakvv4IK4Qum2nSEw6dbGZ9QNyY2SCoZAZSf9auOk4k
KKN/W8YaomfJUViKKkbAm/YvUYoLZhmNtvV3v20ZMcvd7cQynkqlXYULMxhz5rOK
/BXHPBtYpfS+5BoaGE8ENx+FG9DR09dREa2gUWItm+wZ0RB5hxTQMZwF+m9jhCyc
al7jA765OhtsZYVcSMrrs5lpCGcfkN1vzhlvI804UOeqb+B79h4u6teyeGFdRfeE
gL0bwp9g4MYVIwNEp3/5zprSj9mHrXWfNqjQmN2V650VrdnLHM1zQPAGA0+8EfoL
Knd4YTqRNJpSpvJaq2jBdSW10F1OzDuYsZX54LaPnNc6SIxSKKcMh3MG6i8GAYFi
KXSrcESzuo3KhIor3hnj8kNcdWM3E54ALjrrCa3+zBCL4VzzS1W1I2dPi26i4/AW
6bnSjbCRryYZuvsxAcjBTbJF66YmfO+FTNHBtOLUbm5D1wSfQbsw4wBewO4waLzN
csnESe2cwzP309lJEMP44qRIlCRIfmzK7ik82+Yc4VQ4SuOFCF1DR4txv3Cq1dVu
FxbPdDu/wzrGy2+NSMaRddnk/VYhFFktjxwpL3v4hEhs6FL7X2CQ1Z/UgSsqfove
Nk3RGF/IoNrzwE6MNDtYyM54BATggFsW0kgBxrPQohgQ4s5MODQD+QuA+lVauPf/
nCjTtJG+BtkKGq5USq7lMTCyTQA4qEuaRmuFVuU/5WypC5ezoxOISQvrIZhZD5jP
7+N99U3eaU9oJOzGVM4QnlGyM97ny09zCihTfhRMoH5nxVGerTosXWAMHmHIMzoJ
iXaBoTIrFsFsuMxQOlNi3jTuhIWYGX8DhHnQCLC3dUFvMUqJ0Efra9IjLhzeSjBw
+3y7Kkt4daUPhjIpP0TEEBi9u8o1mjXPe1Ewr0c0CJscpfJWnwKwo/OXxI8kGVOK
iM/xfs+mdDpnPARSAIg7jOZ59vWUJ+wpxvYLz6niOLgHWeaJo3s/n0a7/VttcHVG
P7zuyNvUGJ195RZ8QEF/UqNj5krutXWV0aIAbC3B6qrJS6UTsWEuGaMrGH51GiNr
9luFwKDpr+XhGh5z9mXIvNjI/k3a6g/a65dOPKYriDSDlyWNVvTqt39mYytpf+Ih
FTTc98rS7frU52A2NqPU4l+hwK46o+6Sr50HT9zMhtNU/ShA3TTH8VhZja05IsG0
710BNVb/vJMK9CIXo1yYTexif3Gf70/SjyC6t4c9CSmNrVcpSK365C7ulHB1ZeP/
VBlPbYZu2nc4aEKSUCLF8kGUQjt3bzuYuwWMVSoIQ/JV7NbOGdV7D+3vTudLEiwk
/vKNv3My3vkYtaQ+Se1PgPyl/aO7sA3yxoS+d/DrW+uvosuqVXj82VViUttLaNbf
mrKu+wdBfST8vhKiqKNEiYkoX7nspMTJAw/id09iaXw4mt2RwUaxH9zm+kGHQtyj
orngY8paZzXMZeno1A0wNhspOjRA3j6zlKzTfbP+J7TUDIZckrXua3UH4LlmvJAE
lTovbAMdCtWpHXalzV+QrceNDvVBHoYAYBZFjwqjAdciLyshuvmpZHp3qKSIdT1p
D9hIwpSk1e0gA+YSYTgrtv66ZLFXYZQZSM+J9AOV180FwCAMJlp+qiP7lTA7SVRV
dbKXpC4034T3Fs1GE7LSjjoN7qXFvxx/OYRrco4xdcawTG6SbTYoxnB27C4ITZoZ
N8qN824Oa/kSYkSPUoeftcujAHmuv1y7qsnjr7ZFR9ZZVl9jeqoshpcxola6CKHq
fdBx2bPJ+B2rW6bMRLCbROYSEPwIFqBk3nOrtML7MjDAlXIlgXnfGBhfPXuyU0Rf
XY5L2WCFXjoKxZ9/9xSEO2kAMr33ZSCat+ZtGzYqYQltdrVPc9nu8bmyUZ4VQBS8
AiCAnALNbEWF2vDYU5vQb6fG8uxx0n+1xM9M1Kn/nO01gp0KL8p4ngyrOiM5Q1eH
FF13fX/MqI09tvqHV/KugCVe82ypsX7QCNEJGiqMra3OCjdwluYb03aqdITvBLN8
cf9pdjhurEaht2EZpboTv/JXqplrNFNWOfJ3cn8qNG5N+4LsUU41xQhRlGn+UmyJ
MxoYt2pZceYIPzW3qUyDeEFcW7UgWTIULnWrjCeSmBhR5e+19w6nhH9zLDnV24yA
v8wN415dc8ZSTxYY9PL6k4FT0JOh1ywgWqxikXWQQNrS89UN2A0DGYDpQJNW+tyh
3rliHMTngaiEAFUtwJWFjTHsdk3jYX2+QvVzxDF/73240XfQjh4QwPYSXR9Qko37
CkF8gv964voW6hSD0ecRgF2M9hfCBBoazOl2JKWNiPh5O1FJIMSlrhRhz/5hajgN
0dXyYwX4DyF8K/WohiFM1Me7RXLPYVZ4Y7hWgjw/vxPB582Tiu5dhzGoNcqom3Rx
tWw5E0t2/HneSuG1qzQwd3/4hfl3eLhJYpbp4Ni5bYqiqvEehQSxeCJuECbG5w+M
FnDDdc6oJl2KqHqQLdAw59F83sy/H4a9WAJbEp3S37JGf5GFg22Qzr3cZe2irhFH
Q75StCR+lEAnIg5GXEsKsH4Zk8o/fI3WjwmwJhsSpBFxIQg4vPAu5Wg6RkQM0Bmy
R7tI3KLgJhqRtvW6BMLUb4GVeHGJ2oigC1An0U3GTy1tH+8HOWjLg5Yjfn9Orik2
VgDOVHN3SQNX4kRbhWbsHZJaKog25IzfNgNql6CgtnnFYGcRZF8sW4m6SAe3AUFP
EPXmXY5RrKqHN9fT9L2xOThAztvFXjh5sNru0X/A8DY6T/btjgRjCOGCswyygCWi
kNhjo9xBqm4GVSrhIj60ek07txRWTramKIZys7orDCVlrhVhW1CTVDsT2SIY4PlD
muwLjjDwy29rsWoVRvHUVBdx+CDtsExLr3u1GZRvG7kIeH3D9WeVGbmdlyp8KI+9
4IFU39Q8pVZe1UKEQa5crX8EjFPgajBwsgY+VtGmj9f49hmDaHM7Tk4tngklte1l
uBp9L6L4pSB5A8FtzNrG0pQUqUMNsyu46Z4lvKZTks2TTLSF4pNOK2NwxQ1l+Tzs
fa+SDPDgAZkiZ2bLqWHeAK4LMi8YeE4UgPF5vQ3flIBDMu3GFb/wTRvqaHfDV47x
fEoWCLqBknk9YajGAq/0HuaKHOHhYTkpU0cpglDTre8MTAuKSOnP5hANlNVa3qoX
3fMbwFp1qbFephYnOEfhwbRODRzvxF2qdbFQpgccBzyrlM+gAiaTLDt5UNIU3zV6
iHfG8NRv7U/+pkQsNFFeA3SQAoBbRG0JNKtqKbVd927XMfeNZshtaUGwVh4MRWau
PsyIvE4iNaMpmJvBakmBqUjLNhKOUEeY1GelKV5VYOXdUEgYt3RZoRiQtaMH2rkk
I/PAfjrfczi/ze0r7fZmhqFGmmA9qxSZOZbmwSC1OfYtpJOf2BX4qEYTTcrUTQjC
p1gmeBmNQdhW8hgaYo9rfO3mtwzhFaQdYHsGkTm3J5Jg8vtKSg5sM8glIwFprXt6
p1wI3x+nFL7wmqCMU+Tp2R/L1wPYNmDRMl3xc6VFeDdZmOkjxBkaFd1NAbMDYgTi
QSNW/8LksK8jidq6Ib+bpiIeyqEAPWK9SYYh4hRsIOySmg6FAn1/UHVu2iaA8fCh
RQNYhtqpOtxqCLgKuI0Aa1ozELUn/0F1fVaN3PGFFLRFN+9zFW1cEhh+e97tUHBk
Xk4AX8NsVkw0XF4UaYJb0zEffVOJhjoECU7NvIRaUIRBgjUASzNcL3tpfKnDb+ej
G065803f4C3zBZDtrr6TQQhGy+adVaffPZWWNOPBNO8O8YnYKAURNspbxGtXB8cB
0FG1/x38m677GS20M0y6vLB0B2QeY++WARUcCLDWKNueIG63M93WcceS3UwJSw8Y
3SpJtLhivp8WeBJ8WaAUULqdAST87T9RCafIhGET1LK8WHF+bk0NVxBEv8VElwCV
8+VgOJjfdd/jShKBKBCavLmlD5iS9S8IrOgg0TJ8kr0g8aLW2sQ4djrIXpV+oBm7
ezfZQ6vk7+r9RYhEIivC8KKi9AJnlS8DTjx/Kc8o4aJAlgMI9+l4WFv1drynVJlB
hyUFNozPXAyt0kzzica+xd1a11dr8gnwSsTYn9rEXQNk4WpFZTyP2K2HMIYROPUK
doQeOiUCdt5rZ/qgFDctLiAR4GzcE+BxGe7453d5NrWCMQGZw9jkZXz8A9DPl+4r
dlwUrlNesTnFMObjUB1VBToskxnHy4uTmbxBAgWb5MSGMaEdv1Tu/I2Qkd39gAop
FAK8AZTdVZHVRkhufvk7jBQxYEcTfvggTTMEXfnDE9Zg+VmhuFPCQkQqp8DYZ9Uo
q7Zh//PA8fPtvH9f/+hFyrz820l+znUO8uZRboK4CGVh6t9cPjUwLh0HTx/ex3kv
5eov8js2PzLA6LExqZXy0NwKyIbQVQJnMvJ2su1lbEVKT0LByr+py6PZM54o9Odu
Tb37i05os/z98D1KhIyZn48Df0KS/Ds1wMCmnPKEf33ED35TT+z9CINPZOU3m6ph
ChUwEDIe0rU4Uc8kWwzuvD9TwvY3hLnol5f8ykpIu9M03Thqv0PCnv5Hmw+IowRg
BkYVSlciN5+L3exO1eouVaL06GgA72g7z2LE/DJtMunbVmJrDDCxZLzPnS86MUgn
6jpeQsAnBLoW5n1a02LkHSxmz8L3i9Z691Zs0rMVk6OaEbhje5aVUDOfLi8RRYt3
E7VdT13sebErJrjenIdHp5EqCM+8whC2jVpb9S6LQ3uBnseqvd3b2wKL9bICV+do
AHPiiAu0qTRMfvKC2mNZjR97mq+TqkUcBEu601Lu/P7AuVikfuxz0gwFVKAyLECs
lOytf4deL1FnU9ZwztZp99O9rsBykrKGV60l7HZUiAeImSaIje4wfsKwrY+OSGCu
BDfYJNaccm9KyGDd+FRdOukdQVk1wsdh5l73Zql/Lk5jDdcm173VrM4hn3daQq4p
FIK5eKxSvYAylnW872i0Xif0jai6CmKsWbCwqutCfl6S/qluu8R5Rd6a1o7+Og0o
4qjszI9HXCJow3ep5bc8eiXQH+cDKjZ/bKAZ2CuwlWb0dshTQaBT96yKWm7rQY0Y
4nMX3+rc3acSEBMCUbUS0+sJdC4ZfliQ53OL81SmI3HifEjweY5vBve18XvKZ7aj
LTatxYwCitE1mplrDdhQ1G+Vhjy3MPC+5TFgik4tgIvdleJzJ+juKmcw2UnawqO2
HlalflNTM9YF0mOFgUes99/WzOdSD/W85rXPvWZ08GmEWzN097Rvky+r8pysyw1n
ZdA9hl69EcDex4I690pIGAPbWyFKmsnap0fM9HURxeqR0gXF5V+bDFc4JqMWRfUt
yr0Dw+kGDl2OfyxWmMtARS1MF3OAsAN856jZgIudQk8KKTCavVHDP8/vuvg1ESb0
ij8b2286P8O2To4KH9NwWlrKsjIiG4yDGZLYs5UTX3qCpUPkT/44qjkCAKhGWar1
5c2vFuAOfVYWPhcitL/hAnhBJpD9xw8iyxsmYJrS0iFMqG5Y0hRNqIjGv5DlrmFO
gSznUe+W6UmqilxutZsu7pwEoUHPvS/vuPQcv73D+IKnCgLhKeXL5l6/89JBPOtu
QjuTpYMqyCje9OR53V4kmB/8aCC7VzRM+8hqEPzB4WifK03qGs+CU1pxGEMYOU2h
7a1y58kb+i96qYmWnEYVyT/cpvml3n+KgKoy/eBHTJaKWmo24qFtRiI/xdYUiMqU
++rSQ3t+LHX9U8PQa1PF7roxulmUS/S4dAvTBNoAfeLTfBhdF3mEUnAyvPFJ6GpO
nhTynE7tZmMm+F4KKWs9h7s0VKrphlnp7Da71a3539iNLKG+pbgYoFDcD/mvnv3E
zGN7D5sdVF5RrvHIQIitqciwN5Z51Tw/I0teUgJ4jXdbAMSZfZcAYcPNFCdkvP74
e1WE3DxkgdEY+wz5lGZ5+rEChnLFtte+Ok4EgD9dgW4PRx1xtVjtbYzFR8GUjY/i
hu+YYl7ly7GLe6J2Yvch0BEdnzVJXH0DT/wRAAInmK0k2g3GnCWk0Crlv+FdUAl+
dqIsildmCVKQv+uOp/Qt6qJBzW86xdOd/YRXmO1E2JnflBO6WBemEC0OpI1+wk3O
J6u8c8m8CO0Oc+ZDjLQ0b/uiYdHOvXFhAT93UmtOBzsUO5pBw1tAay5kBth8VBRE
BWfNDYh7E7aSPwf2nO0NSyEdTUoLs/pt4MCbD225knmFFh0jHVa9iRgj0AB3bttP
YJilVOFEgP0oid7Wd1HVaKBoMvOvmNxJYhO1HffPbKkQI8tdsdKDUhqhmBSx9Kdd
fhWAAil3ZFdgPVfJy+mF4NzyHouwZ2Nt9Lfb7R+gJsVxM/ZTrTwApgRJefWvnQs7
16xnwa6oFP0A9pSlFMZ+2GNVVY3PWwSRVMdjgIyD8utEqNdnzD4by6BaDssMZmtz
aDsA36OJ73JVWZilwRAIS6LTLxW9zn1D0VSyYdjuyRAZ6qN2Dw/E/Tb1tUH/rP56
yoeu4qMtq6XhyhD5a7HpoJKZA1H9dqprgoDMB8tGeLRJtlH1MzAx1ha05701PpRo
9TtkV69q31HRFifjXkdCS5HPs3bg7/i5vJ7S8zQiRlW7DqMTGUpCc+rRtVu9Lt/0
DFw0q2itb5Y7ieYEic2iKtM11uDxrQjlUkMvcYFeSd6Gi0oT6fi+OX+Phs50uNai
83+PrJCIU8gbPAeUBNkTwFBdtyjORmxnVDOkCrHPW9M3FQRgVQINQEypjd4oy7o0
xspXQBvklusVFeGcStRvjZt6JpzmEf81gKcDv73Z0El/u4AHv6drlip0T36c1Ljh
8Xt3hcM4vMisNQNCMDdYBzOmh8ihqR5JZ0GhxjS/ruH/roIiMEGjZq6lTSKkzq+t
waggyTa/8ubLef3FRCA/e/pQZF5PWz4xlnNDB9yAVbAI0w3Xait27jT0aIMNJ717
Kb7l88gF1QtaJq/zYKjnpcECuRe0b3A75MiwK4fXM5z6NyqRe69jSeL51nWtjT5M
ao/VJxMVaAWh74F4b+bPoNIjZdRPImRAbpqW9vL13MFXrdVVtRO22IjdeXmXxH9q
htyQSmAhnMmxmojL0C20x6JYm6mVjjxajDE6aPAVf2C9oolxFL82A+QTLd/HUgIz
gC9Kl14AwHb560n54ZCVeMl3J1JIpEEVsV9lEC6h+7GJB+bZQGi/kXzPxKRN+clQ
gdhXEsII9vMFkww9iwo5uh9hbuZ7O0DbGiWJcJTWlyBXAqkSuG0h/Z5waZUHEUjt
t8b0bV0IBkA9HxknvJ6RWM/reJEsU8zrwagtSx5t0fhaVTy/JsvcsevTBdWb3ChM
sD745Y714l0q+POKzD+QdsN5KhmXF8u7X1IvGUOvqyU2rO0gxZxxN0GgIqbORnV2
NVkJXbgnSJqiXL59VcVzNgjyvqk7VhQmS5DQOSiV5HYmY4wV16uwgmZB0CKU6ETM
5tJMoPYSrxtXZgtz0KV90VWwllOn/KTT+B8npC8Mm7JHQjMcUklZorHxIyceTBw2
cVTOSaRdxwfPxrujVnrjUhQA7LxIBsBWJoVAgnlVSPCw14WqkOpjOWHW4gGXVG/E
t8HpCUKCsW+FbRlejXYHU7B1dKUcVMp8C0/8NG0/juOJwySg+UaM+N4eznbN7JRy
U3aPjGaPxbKi2osUhfvWrobt7cBcI+5ONRYkH/tKb4Q+D59BKeeRN9vnhkqq3+mk
PcFxW8QeuCza9Ax4K8L92axmkeYTmogBFmITP9rOB1b+KAs0CV2SkzSvqOrLuNlh
3qG1WQzIbkWxMrtxM1EI7qrTq8zHEW1fJxBlNgkP5n7gf9rx+c+sGi5t4QvFF7DN
OnOgoYsdKB+A4u3nMxbF3x4VfHalPjGvjoBLRiH2/ApOI+7OiZD7hkQtQJZ+zsbf
1uR/Yx++ipFVgrKf/xGgPMhIQ2SeEJlzMbWMs3kGtVeg8L+lr/jr923KjjIX1FtI
0b1NErsH8qmcZBL2W7BzUkIXr41cIngNuv6rFXdQaFd566WVOy4JZdlvaWRPSAqS
1+WQHEUY+Oxg6V/21uFdERFte5OL+dEwUPOeCrlwkGIzI1qgS5wQLKcUt2l5k2ES
xUbriVXEQjnVe1GuAdZzjEXLzrRePsQ9ThkQ/187st+Bmltx2Ho+Ba4Vrc2jn+FP
xvA8650ymVKRo0C2pQom2f+dyk8bgCC1mF8QBN3eAo7GxK2sFR0VXal735iZQwMB
FiHPq1KYrifFbqC5lrK6SWZ+V/hUc52wFeLI81MPiKY5NTVUCLP7V/B0I+VW2U04
Mat0p9tBaNRVR8u7LtByqoFT4hc/nKNDIoSdrZfpUPylRuaKK00EivEMeXigzZNa
gyAVa5O5A1YzkjZT/5Bpm4s4JsEU6U4Zl0sYPtg+n2UtIi7MMtYfKZb7lOQb2Elm
p2gBBza+kzqVYES286vm5Hdz54pZAVQ3Jjqw6mQZq6UFKpwFO3caC2BehyQCzvgs
LWLiXJn+E6SdU1O2KoZwdkLJIEYWT/1V+bpQ4D+QsJPsRZ+b8ulc98M2Mp0gnlBG
VriHHqHK2ZnJx8dOS7ukspDLDXfqmxEcQ76E6JxIcfnIHkCpCpmqH2sPknt2p9rY
Sm9wz9mnMdLhXcBRiE0HXkVbvZCBUNT58UFesnzyGnv9L9VmoWxzqi07usYSHQPj
+cZcXsLEKT9pvpvnxnVL7+H0WEHx56qeSXkIEXgNDcY01pgJXwHTb2mraMU+dQiy
L8ipOLRC/ETkQVAyWR5l11Z7dICsjyb3/gxoig2T4ZLKBg1FW07knrbbT4vqmJ7Z
Gbx0lAWzQjaGHjATmNa3sRMvATn9zlzeXOjBn3+BdN1mKuofHM9IYYbbI2mufFMz
1WQ8qlPmkqsCFxZHNWeUO+7MoUmfgl729gqbpo8m3C4i6J2jR4T1JbAG/V6mvdT+
WL52qsOruiVxrtMc+3KeLfLFg/SQUtTaGQVVspinR+7Op2FBrrT2kXP3yKV03qg5
FxFBBij1omTst4+ll4FKIQwOb55rI5nH6Jk6x7aaGNiFz85m20uofDytGBJWYJ5/
NswEgLFppmqpVlFXriECgwDOFAqjSs77zTCmM8WcgskBqCJlWwomBJf/OtJlJAwv
Hm8GX0ZDq3kHDHBrButxqDjb+UOzQJ0ldcnni5DcZbbCqQtEoFeGc0lr5CjEqTtf
nIlFZXt8Wnn+b8g05kNavzeew41d6UniPeULe3YyvcvlmUyXvU3zZPFa/jaEc5fG
qae3RJ/Ej4DMOuugfFXsHcyQtmAgYannJxPs62QLNF8TkpsNaGwQbpbwlv6lzHCn
Xx+zIbu6UG01cApPeWOZV6dG4xC/vzWkxnthkA4DcSeINV7icXExBmJzUreaQCuJ
Q/fJZiZb0yI8qkFgi3h3F457PfJTDKSZ/tkUhFBmBvYQ9Ek6EzVw9191kUjooXyM
Y5naEhp5wjWuMjb9OfUKYxmCZToWlnBcGQD45PvdpoBZwrub0O090Mg27btBbt51
nRa/LkoipgWou94qyO1nROFfMVYMxRQ6seQ8C6kmDP7S7uOq0iecDDCa4D3JIp6G
UC7RGJX7cdWswswOGnE3CvReS0yBo0j7DjhtDPopkCcbJ1h06BbjxQBsHQCevsgH
qaHmNc2or4wMPGVS+jC60Jq/hdoUf/lJApX7nfkgPwwi2U0tOQt3a+Zl8G576T+K
vU8pR27yvSLowsMMgMOaaopUkd6ruqRMAilHi6j74AkpHROM4HmeELPSldhoHLh2
g5LVa97OB6dNwh3nEnzOUhliWtBo0NyMsyvLPKskeuKkGB1H1tqH/YWFLeBGqJ3u
PUuE68H30W9ThdbtYxaE3I2T8eHAQ5WW5XA4i0OeHNjuaMBW938SMAzintKs59ek
rbr0tmE05cP0PuSXj2OUQprGam1kjuiRr18vZB1TtKoB6ckrcxp9uljuZeFj9jS0
87HWLAF1Ba5R6r62W6v8+m2ge1fPRVr5kTcHwIPgGdcBzBdBgEh/3+xuVXk2e1L+
SOFxNt+2P+5BlJN4J8UfQwui++z8WcciAzgyJJGzrRNJoe0jvvSnKIGQfOm8LHyt
MVsDOQukvZ1zMh2gMOTZqw0IjJ6J5AdChp0BEr7vMHR9xJwjhYtNDl0EtP9ZNGpq
5EAPS5kbxvYeQLiTXaExjwQj9IgiWiadO+cYWYrpcnvA3j8PhpL1pP8P4umO2X/Y
t27jYp71yGbQf+PMIdN2WBCeL/wawRAK4zPAwh3w/vAcWFK54DeoXLYmYXX67ZVg
XrM0zfHH/817VHlCnuvyvTJ7GaSkU4mLPJxkxANcVnhScafabx9GTdQczOXoNSh6
cHpC1oOp4Ma7I3d+xAkppksmGMRcC2+xeakPm2lZdFioK6YlRe/YgKj7nAIlLLa4
DIwSVgMEXzcj8C1IESxJMYJfj+zs6XKlx8Sqdf3Bl9EH3x6UExobiqMzAe/zgrEq
6BG/kRNvv/hNomDavyPmoVa8Iy9NBTPs1z3lsOzP54p3gneUpPTUYjKRuJWsm66P
hDOlGXJanIwA24Fs3oTnrnyU7PcVyoWU8WBorRIoG81beBjLC6b6NfmJrgymydCf
JBAq3OyTgHfb1CYM+bx/AWxHldukDDiPsRkKQcE7MGQmBZZ4eU8jWB93hPxZzgYn
RL6i4fHKgxopfDgDHUechky/vI3wuMMx26q1PWsdim3f6vZZryLQ6DQVZZC3c1Sk
UkWBvdpkNY7GyG9CSIw5pAknpgslnVhYd05Np3HnS2hLwEevfo78thRiZxh5qS+y
CZt/+sjl/nM3ozEBMUDYNM3UBeG0UVReuIMkTADXEvG/EinLO5GrT9ZElpz3tv0Z
mAbTJMlkjkVaRwCPTxAS4WD0PjE7f9Oa6QsjCHbsdg3ju6akXQOMyNUX1mLWunxK
jmOw5sRBt+RpGYLB7BvK7vUHJfL/s0JMcS5n0vMNM4/kR+3UXiVdJOWMJmxytNlN
ZJ9inRI7ZvuOjIIo8W30TuLBcGC+2s/5dNYikQn8q6LOj/SUa4ICX1FyiAHfbzVH
IRhkrrOKxQMvNUvXfSDI3pSLNIPd9PwkQqc9bSGvHKWosGjjKTXL/0wcM5NwhBVY
jp9/fJdVyI3Jg5MVIgJWehCkFvy4ZlA9qFTrkbw8I/XfWsT7+IO8UEZqxsTGhAI0
a0a0u/eoxwxCgSWnlZIgXrUpSFiW7dXRVI0yuQHEEGEp6Ju0zAhlAtp2IxzJkaNj
rI4uLimZaTzEV3Mun00P0JPWCxj58ZcP3d3aicHs85PIdQfcCyVo/GCPEbvDzd6s
2DK+UTzOBB0qqYcMKXuU1/YOGql8bDmF9p0jGFQ5eMe/hHrPevr5WjmroObtXIDT
nCVst0YMsE5C2iuabRoAXz+ZK6NU1bSe6KL+Sd2mMrj0QRwZfGddBU1XQEj3xDWb
hyQojgHSLF57NybGUMdMHaWA3LKq1o/vL+C19eurqY60Swte1yrFjABJgtAo+Fud
MM+kJyn8FboX9BvjwK0oNN0JO6eY6ke5qJVW2o2Z9TSt5hG+1xyLLlYah8Y4qqeR
GdriyIS6VoT6Fh3jAkiQ2AsBkDQ1UUPdvYoR6efMkrDWJpqb7vCwgGCbwl1VJtvl
4nivsMjF+V4jEEGaZCvRneOqQrL8yZcjYH3Srevuxm8jjiupDZRumqotSuAGurye
xFNjRVegshwOfqvVNPx0iR/r9qTKgfjnJf+smpBJKUkowhA6svIOUguEIaJKGLFC
p3EnB0IjzhKhlRiEReRhtUWGjTUPiix23EXcu1l46gHuO2G7bQSyH3rT9d4PUKQT
Ejx9kzGAOdgf/2LxIrgqs/1p1Hp5sweCx5CEALkHoB6oMM6tzVzVGA7NiXLR79ly
+jlknUWwHUGHycSfonGM+dsfUAA+v+lWr2ZI2hiXitoua9WmKmLVd01HKJBIsvbQ
PKykx80UXxPgMr2yC1bvdZki3PPy/W3I4NBQjai/lshWeW3dbcDwEgzvo5WTNgQa
QkovIgP1Y/HsZvcAeCqYLjT28AzUgNQyIZgdK8UhV5SuyrEaU5Y9ZveCqp1BiqDO
o/GbXVqXRjWvN8D0wcXoPB09HFHnsY3OpuhOPnaxj7sg/iLZRqBhNt9kd8UXcFUO
BhNB9z/OMFwsATd4ekVDliqIUsFKghQeLRUP690Mtmxg2ITTxJ1Nv5TuaImGSZC+
IXHfLBzOccYNkfHX/hfOOX3XDmGF/tR2QoXOycIfsqAjjdNKp+Dy4RXiNptWCGAa
yANA2dLuYU289eDMHGZxZFGcd1i7R4SmstRixA6gpSXYbAv2/Bel3UhRFaN0Xpey
8gnxjL0FZnMi6JvBLCMqalMxPaRYa9sIOECoAyChM4LWXg3fVbgmbdN9jsPaR+87
FSHQyYmGBFFz20GexyYNl7ix2YyI1y2CM2QjtEYbS1N6U6HHObITZGYh12rqvP8W
nSkdNaQBVGwMnv092AA+QkyfAOVPbhqFITH0DCJcCQUDQiAcWECW0pjYAbfmLq21
c0+91OlxxdiMQW97qqKS8ANawtzz0pVuSKf+RRwoXfpjWoaCwjbW/q1JOqMryI9x
HKqHygdMb4hEriIJxwTK7V9uRYuFfYFormimZJA5S4E0Gq1oNvzbvO+zu0TdUtEn
8NCexJLoHro57OnhTnhiubfCrDGirxqCofhW4dg7FTXMUj8c0d+CO4xEdXA5I/QM
1sSu7ghh9qz07O73pZFTpf8j8cGqVJ5XaKwejQfr59SVqZnRwDhUQVxNQ2jnB6Ls
yeSX3ZblE1bRE7n3kMckWrluiNjmxqxkQY3Wb4nTLq4vN3As0lPMkFSsbdZcLLRZ
Lpu1Ki7StLsAAFca1Z0CEhEvnb7S3cC72rvtC3yUCob1r5MLL2mtbzF+vu26N9lg
jZ5oR7AGs4yjx64mxteyPVWPVg+PxTbMIVdo3lpIUvxuw37Asf2Vhg7kWM7+nffJ
yYRNElfrFhdhcKYDc2HopgVxC/nZ4bVVdIegYjVkoxzbCUuCV1vTv+eKKOK7XkEz
qz7sJgQHVFp65cUV/UpFEIzGYQJHO9OUOCsmVAnCVTmFPSQ4cwkbStisoAaAil9K
ZGo4PHj5MhuIRZ3W6kwbADnMV6JN9hJER4c9cdT2VQpGeY1+bSflmhhPpVGUQhfg
+BHjz2t1W0IqOp9q7FaBzhgMLXXyrgslryU6nuY3SvrJqsENi/yZnuiYGlhPuP0x
ptaSopzxuLrnKcnaNvcV327szPXS7hUqeD+ntEWX6ShAR22ONL6XpiGOpxJtCj8l
cARoD2P9KLxCF7f2yPMnIjpIi1cisC5UZp9dReGZA+lR/YVtHEB0G2C6zE2wWreN
NNnALoMdJEkBVVf402XdOkVI+BSlyazeqzTW2d7qZrItYq70iPcTkQyvrv/trorx
50966N+1CnAjk0G72EqLD96SRB94x4NJoF6NOkPdGR6Z9rZ9gRuPtnoaEImeBkHF
kpPlkDDV8JobH7JB/hmXc0ScaoXRAAoKNew1e90sBe1HQeIVb7sbDggusg7uaMqt
YjVOCTOsNbflx41Q/6UZVMc4zOJM8R4BSgvrJ8uCO6YjS7DQsl76bgnvakE1vjCe
EowgNxJj27rh0ryGCAZTvQsGtv4GmeEWPzKQiVZ7qf+gzSxHez9nfkRI3NMwYRH/
MmyzVSI2CfRVhWd/y6f6oVaPPrVc7/ZHRZ9gox6ue/QkjHLTuWyKwauzvxPeUsK1
4wuZnf4B55bQtxQd9wofdoiZz/DNoa1bLEf6YBa9jUMh+OVm7BlWFj47WN7TLfN7
wSJR7qR8v62ma+U99h3q9AbX7ajtOGfyHBsTKvp7nV7RMZj8AguwWJBX+lHzWADZ
NPy5DOOMbBeB2RG1Mv6n4zqNqddalFDRHUUwZ9dnz7zkH8DOqMf9lrFfW0WEztNG
GSEDaKSCy1AYpUVJIhTjZsg/95ngPd+f2USiv1MPt+NOW0ZqKA3J0Af+IUTW6IeO
NbiXuNT+7C8pV9uhABpvOhG2MzRZY4U6BSj1B/cjofUgguZf/0eIkrFt3A4uV3DF
2FdiqgQBaElX+zayOeBWnqPc7A+BppI66bBoDySeJHzXN3ugdJBRSwxpzq2/e6Je
AwznNfR7VH3anHCb7aqODDQLUMoNilyc5kpJrVoqOyOpsa3v+ybE/csdz86t7SsC
umKdoc+nN8LMdtRbE+nhDJ05Uqh97Wk8+IQpe1kkwW/XAWhDo7GzngKCyYukXEoU
RJ2QNM1/0nKx79y3qLgfnbSmrUHuEOYYbGsNx1/pbKQhMjzs3rSstUV8wvMbBN0G
93vOo9ME31naAuL++kUOIbRlBwdZUveB4pt0NOMV/9DO0weBmqIlAdrQjoj22Vfv
JWhOZbvXuCEYPITHRbsl4yJwt1OrJrOSjh3ZK6MIkt5CSJS0X6fucj3gkp013kwi
xRPnoAWXrkP0D89Y76jjxj7NWYWkLlWYX5yx4bAx2Fp5+fQ+GgA7D13fHLfH/MRM
OpLTvSxh4g2TZyfQuPpax6omiLNQ//j3Yp4dHiGkkWPBhiI7fm4GM3ktyfO/28BO
7nDtn4zVa/pIVcvROLmaWBqhI8MViE4Dv7AwG79UFPoLPlT6q2JFQwE+bC7IT7IS
cLHSTF1n2e//5khqVCj4A5rqJev42OOGS3xoMp2xNaDBJBMrShybgR8Anv1oYz9V
EnPartJ+ruoXfXNtGmy/GTsIjX1IFsNMINpVx6So50JNt/y2/2Wpv9mMatadPfaU
Jk1eLCjo5CpXuf4DOuW4Etc9pebfnOrmMiwbT01yJz0xb7OaRccuneYZhbR0emM7
CVMzF4MVxV6ltcTjnxlDULERLSpB+nOtkWilXFtyt5S+the/B97Fk/Qj0ENdyWs6
QQGB+NMknSNQi0FbjRk1dRvlof1QnlIpgrBDuKf8sIxm4ee3bdH9Cse6SOSt1n8Q
DGGIJSL29k/C6Yc+4tkdgC3PYn4l378j/ksBBFDBB2dhiI6pgJUoNK4KkXYX2WDy
fZlB5hpIXo/2fAh5ZyQxLi78LGoxXUNRdJQhGehk7O6MKzYzsRmG0NvuAK2p8EBx
EmsT61Qg7Wryaxr5s5xNCzKav8anAfma9Ius9YMdqlYsgJZLVDsvsK/L4mDLf4G2
SJlfr2RfNfMADtp3uLXjL+A/Hi2koHa9wbTqF5kDRWAKs0AY6hzMXOz+F0G3QKxr
v/rLgc7Ot2UhDYO0nXLt+IWy8PGg77Et+kHN0uSK2p9MdpVPHyusA3kJGhYmAdr5
5Rnnl+1UMBZz1vxnlKwAu4iDr1foOtUcu0GaCe/dMMeH0Adhh7evcjl3DnXaucaV
Dw6bXVWoyGlMb5Ep7NMrGYafi4tTD/1DUTTQ9yuk/Fd5u7Zmt3+80a4zm4YhSwNM
JHU27yrmAQK75SeSPqNW0IoeMUTBmH6SPwf+0Oe5dmVAadT3FpvFv+IjuF1WcSB2
sxK3IN4DOWLwyT/r4IN6suT8Wj5eYu6kZC83Xao+4lkdRwcI8zl1o7O2eOWRYsb2
K31OCzQNDS2681xw7duJ0AU0YDP+1MZK0yTrP+jTBVQ0wXUGMb5h629DZG97fAXa
U7oGXnhawwiq1jCYsDBsU+Dqdlfj4QfM+fE9m59ydZnbHU9LZ9p9Pfgcu8EGgZfn
j7TXZRz4pN+TSGt2yNFWD22j53M9HyoqsvLyJQy0f4yYF+BRk7K0xsud/VingnPY
KOz/N5bDaaCzWNRhttGkye4ubyfdAk/H246pU87T4ZHZ4ZXkml2xJpl/HuvpB6+a
jfPKdEyu3/msus6glLt2gpsMHIZcFkgG4DWoLIKIy36iOt80WaOdpXKyBxiNjdcp
cOXqXGkrbvgE+NFhcitAXdxxiFbi0GfKneJeH1wcZPHNq4j6gRV4/ZxavNaRN+iI
usDLl8rlaJ+cc+GbPqvfxBEqfK7E3oCJ1WAx4tADg/wVcUSpkPOF+DXQLpvAmMmb
3lv5yFf0YCaaMpsOn5ngGWBtbUc4fmIw7jAGgodUiHrDPDoGMmSOYD0hcIYp1oVS
QCfbtwu/0cimu8J1JIcRs+9gA6fRzhn+eJa3orrsSt1oS6G5HLLJaLFvqmfQL8ks
iPBpFwLP4CrUGLjb7amuYXAdAbq4mVKY5e6T6EKwPyYaTKeDSHteMBW9FWsrp32s
IBZEMUsEzlqMMF4rG9pvRzc2OzD2TSb34SaEYW7aTk6ms2yBqRoc1I4HYZTojCcG
yti2zBwM8TeVDdIo6jMaorQOI2fmOHETJvSb93yT/4E5AD+hF5TzIOGh1L5POVZv
+wHOkwgeOW9gma3hg9Q1LwTJvGCmhp7wbF8zlxTexIh+DhYylkfll9M/uiIYMcuZ
EMoDGYMjo6tgMNPT+9dCw+2+JVHsg3BZzy+h8RctujaA/vsaOYd13Y7rQW/ERcRE
6DS2ZgoCiDcpZIS+nCLB+mNSJdc+KHtdFtkve6jubA8YNQT3MZQz4ZwYr20QsObc
FMuAmElUN7eCYgIr5Z8K2YcG8mN7IjxLgH1ZjkW6YSKpZNJoz9ds6C0vatea2zCo
sDPus1lqWauYIQVi2xAF6lRx9HhsiGo8bA7xh/y5fUZm0vq8uN/YiKQBeIi3Y3H8
CMC5WT7V5Ll3tAYbf9jTXvX3oDxAHWxvNDPpwm7VV8iQ76T9mvv4hOP/AZnZxcoJ
xBVsQooJcMdC+WkEaNvhdHTGzKOMvspYf9rT4FWYWi5rURuEdvQkXaiCDgV0OXOq
c4zcL/2zifriPm9CQjukx0H62CmBfEAxn2d/Dfw7m9fDSEUDq+AU0EA8uPFiUWPR
1AozdYJs7epz9id6GhJu+lKfTcUAGiT2D4vIKmeYJpoPbbxZrHsLK7qIwbAU5sGA
STxRbl2vEpAk5Gx+Kxk9+0xBOiVRZHEGZ4J7KPRsjd6Gfoq22sciVbB3sXMIJKk7
G7ETJxFgVIguCbptMqdnPFU+Dhi1/sQsDB9k1ZYyI3w27eo2t83JQS9c494ycIw3
M+CVhi/V+ZpkQ1wJEDlwXMGYcQ4W5igVjvh1GiQqP6vLvkekLF5UWhkZLrgid025
VBrqh/vRxbwNMetZ7gifpmOyG/WhwVMJfscQQb6QpRIKiXtHcH6FSVu3Uxcdzb2t
zUBsDtz76JHPeY0r3ytu8kOvOYtiW65/+3BHN+U+Luu4OCDsVddlzHggc0bTsoio
OOGnfK60sGlqusha+6Vr0DE8ozCliHnOFFeFP4Gups5AdMpbB5v78i2tehU/WqLQ
m8GJY7ZrGNWHxoFHJK+mQk2dSyGJymteY/+V/boqFPrAkoH/uIBh/ix2Bg5LFkbi
jPUS7rGbRkjFiXV6wwJkWtb3xOy4ErICF3pruO+0HZPjS4KdYo2b+UYJ3UpfHbfy
cfzrDAXqZK1mFOsRZTjO/FKrzn3nen+fXUr9RyqrSYcz7Fc/N5xZvw47zgTP0pWx
r2bl/KvWc9SNdCkgxmbn/3iBWvWEuZu+um82GgRjsf4QP9yWD2XJaH5vtKMwMewv
jRV/1IqeBmZCdgHWJBpL7N92urnZQ/iNe0df7mrWQPRHJSMVLWcK9FRs+oii0a/Y
lVpeRBfQAGW0thUyBrSB+gk0OMUi7DVK3UzHGPk3qzp82AUiUaZL3dL9K9kF/OFk
y2pIR2paf4uvZcXPUnmb+8THiUyMpbmqid3ttcvJQ7ydYWiST/jGvKqrWrCp64rb
dznjYJrwFcb0+B1QXNnyRkavzne5ezDHZt6chX9SiArtcIJKCmmJUNd9YQkAhdpR
ZCjI9skPUx2lV6sE9Y2Mob5wWRSk264pKF/vOeqMtJ697HGGuJHRoJlsREfC5bQp
pFPwXwEr6nrXNDXqwXgEthPma06b3jA5/JvgC5nD5gHkhThUv+UPE/jhPhFg7GAV
LtCXII2FZuM2h+n1aJvvczkZHfUzvleSYv0aDEgxVJghp924eYXi+cdH36fsCxO8
wXGkz5G+Jvm08B1LrxfvzTHs2Gh6G2douGHxacWMjXwSjq7q45DQudDZEnBcjIfx
zYsvMcX+kmivekaFBNGUQ3movyMl9sqhxB7JWaJNuHgwNP2W1TXCuqTrZSODPt0c
cQfGqGTyYAfeKep00DHVBVbWJZl0RyIUVmnBGR7xIGUrhQz768OzGEMD6PM5yECo
NcC3tHqgvEHtNcMofZZAbYRnhZFGPTCK3hNqsog1E03zYA1flozs6ZxnyqQ5rkcU
vAt40OLy2DgT1NeASmgXBSAeRLArpQVMArVB+0DLL0c+NsMo/FXQP1i+Q67I19LZ
aWg1QfcHfSBLNSu8zGzHW3yD9hyfnDZdTeUsXCPh5Z+/nIGJw4nmFsr58LQiS/jc
hC7QasyqGOxVIopVGC9dnxBwiDq0vIyOO/08cFRWCo2F7lDQUdaufvF1uUgArzbd
BDBQc8CO39qQDCdP1U1fW9CWmr4x2YS+A4XW6WHl7cEvxbb8Ekr9aLqE+gwu988X
SzmjZIaRo+nZrjhV6LQLDWZqsopUwKY2bxsEM9x+EfipUQ0+viw+Mjz0CAD0ZK8n
+8CPJ4pBUIom/O9rb7CPbEcSL7PQJf6bfMHGuK99yyN2ZjWfLIV/JIbofamG96lR
guctU+bW5Dy/wvyeBktJDAm1FhhW8vtb0j2hK9LGW3HcIp1D7/dUKctLzEEq9UOa
S7+vtjDyzqT8faGtwgaTRRf2iC+g0KwhEySodnzSZ8arajCVL4lUCTQs4Alff4Mv
HhFyx792hrYNl1JmAlA9fGDcXKrNFEtJAQnAuVgdbX+4WNrKFkVSEVL053tTVBMT
DI3xqJIL/IAeL5hFBwRoVQLABz0HnGryrV5mnwIqHOdaE7Rxn6ljwzzMS1riTx/J
CqYk7tIwiU4BlTbOIJB11IkqnwLwWZLAtM4YXz9Td6cRIXeiC1fvyKfLByC4qhy+
yj1ej6d+3wWFeZxeP+yqQc138t1tSJ3cXsotmI8m7bjN0v5CbEcJ+DK+P5EdMeVm
bX7jrUFNf1E4bClO2ZeKy42AthTDhqvyDVc1pbnO5maKM62/QRw4EUyN8DsOxXzz
pKGtYCQy7aqLBPiBv5QwRUPo8dze1Tw6q2HFMfu2eWCJK7asLUmiLQA4e97odICa
vKm5mKJxQMOixpdIGWqPbeAasiNPcT+g+334A7kWK4KHJq3XOgH1QKSlPbdq+F/U
GHRfqAzpb1fwam/nyphcnYSTfayIYLjl70/XSBd8Y7foQFmGDjonPcuaONPC+qw7
n9Ml5AA7heMireKq++NOw6OVXedme5AxV/j+jNhUYaeIQWei5U0VoqXQrUPXQ5I+
FWH/UP6ptqwG33OB5ypJvjmMxx1IEzHOXmxM6kf6jWEG3nXDFXiID09VIANr3MoW
rBSqlxySZPUJQCJmfV7TSpJM2j3KDA1YtSSffu47ISliGKazH0Omeq+4dFo3emWB
frwxpw2uQLuATO8daolvqphpfQqaNEi0jCx5yNV1edti/y0Aw/9RmGG7n104a8Ur
D+R9wpcgVgIwK/roIB8qNs3SuosEb82SI8HiBXfbIqkuR0xKoxXu3JHgSohkzZ/c
Zo819PRqIALlmWmqPFIoHs4CjlmmOeMAuXIt5oe0CMK+fJ5nATpza3flQIHLn/wP
/Fk10HiAVVTSAva7En0DxCplGUXSGsN9D7UszmVoBy9DW+vCsaStjO/Gs0kbVcO9
bSUQJzhs22jrD7NyFD5CQGHZnx+GV7wS/J/q2IVosJUsJ7a69GRToPNTkLh5Q5yH
+31qn05KHfgOysP3RYAwTgZiF49ImHS5Zs469RP6gHt2eObkeN3rVMsWRSoIy/J4
uixXuPbX/3pSxZUXqfyQEF7fgwoVwHx8ZpKZmZL9Qn/JPSkGAxGVvBIijTaj7mKL
2muS9gGxg8Akj+kxlx2pEw1PTuKd0Nm1yX+PThLQzztyH7DqXAFl69Jj3twjYzzU
t8NhADaXL3+MARjtKkrtMpwszGKPlr04ea8zZD9Z8EaT1UrYb81/Uyt1HKT86Jwd
ylqeL+FylsP0F8WIot0m+qusSZMldtxpwE/kK5ULUcmgWPdJ1dqljSIN3M0nxA9R
WLj3uKoBnwuQRcXp126DdN6Kf2cKAmvwR3voTzEzV2top0L2HvQUFaOqHI9LkoJT
6Tpg193v0X3QYqNcV42a5ncqNlfNB5gr6CXrW//TyNfKBOUdX6y4gAiY/berrAlH
ViQpuExsUn0ES/4wFCvGEDTC6oXy8drefoXs4wPJf1Al4N8OCIePHJ856KYEcsEy
rczQoW8KHwsYrzIMdS1aLs7ZOD6Nrkp05QVWWlpiwGiMpMGX5U6TkrSJdIyjq7WK
ucvYvebE21mojMRsqurKlCPQ1VWPz/FVgsiVUkUaxdNrpFT05j4g3xYzx/bSua2/
8eHFc+iFnthSKyTphKiUE9MCCcN+DArpnxAjIlM5EV8BHjZQFTTES/AgZuu0nshX
FzwmQcLPbARVAvRbHR59vaNG18u5JiSEEyf1xkHdj9PVF7rcTrTYkkupy1lIrY2+
hIdqQHceSCCsvY3fIeZITAIYj15R9XQKgsWDgtgn/iLxZ9/DMAxrmWObgltZ92wi
OndqAv71W4egOHwJvLOx418UMefOyW9//x3yg9YIVPwyQfdsrT+ke9943s0Z9V2Z
G4oJKjt3a3/Qo1/CaXE9fnv1fGA/9XfUnzj2CqrpghlfONxxCnQBAIkaG0XVohmC
2ly0xEO1YuemcjnWCHa5J+n2N6P9u474CK8hTPUBnIdOftKtniyjoCZfUf/JCZkh
T2cAxgLEJAjxtTlC528dNNCn0FL+iBHRL14Fiv0IvFgecz4OgrwoyrZ0MOQZS7B8
sBoBBX6hwMzCOReIG6/+y0FCOq328vBVNcCjtQ1gEP5fDrOYGs2Ao4j2pXxSocX3
YiT2n52NH8tJo48ixuD/7RIdlsqM+gXvSer07L8mizQ7TVfCsqy+bhQA6PuhAHP1
L3NmRtmgd4j1PsJGq/Ao41MEqADOfs1ZkIzMAJ/KX9u7d594BiYG7UyrOCLLTFIT
juucNfcP4Vj4m+wyA9lzyOMs9FL4lLeBlOKBm5euR3lm3BnVGsWpjEk/vPN3eji+
nFScnbBwf6byhqqYAPVYgdxwfa4BLrW8j7QcxKwoGoawxl76I7T+cPL3R8sjvS/Q
LHCVawyQEdeFeS95PHUfmGW0msgYOsr5LzZPyPcrSRQaBWsPXUi5qmm6yOm6jCEJ
n3xvyTBNMyyc4zgD9536IVZ+tiOTjJZkY+Z5AlX3x589Nk+cKbTP1HPl5tUmPOmf
Z4I6ZNmADCGZn9+AAiZpFLNiHMptpjTkmUZhTjUwlyLLp+Alel/FHHZ0hTezFcpH
Kdf0IqX9P+Iamqg/zh4y6e3XCLo5mgE4LqubeSOe0FMX+d1W5pZBTzYsgXp0WsYx
sl7pPIJchqOWNViq5k94AtgM+MHlY5KDa6rZJdD/Yxc1nA0A1cp2lvUuio95c2lI
F9AMtIaExRS8w1ZX+BI2CsJHyS+RRyIB4sQ7hJ5LNgu+ga+SRQxcihRx10ucjoMv
c7sg7sXGEjLCqxb4NRhQXmvO9bG8DQ03YhilwoRawRhRXhJLGOtIwUyfay5HC3+K
+yCB6LCkaaP3nOmveO78Enre0GlXV0Ujcku8wkTwOzbGy6zc+Chu5ycl3S1w3sUk
aqIZwsO+83F1CLlmqkmUWJu4+DjJIlX275eJkzd1aU1IawaGYQ2cwuqoYYJEBkas
lxMmtMTwNSBXpH2yVsxSVwYTNxElyfHKT7cH7sWY405MgHoJ5JuGhtwgwNZj7Q92
rR2N2FPSBXmWOW2yn6aiK/2FCMxkZHoVSZ7uuipfNyKquWEX5qn5U5Ijs2I811Ur
zW3ypLvcYOhFT+wwwK547i4SBk6qLnbDL4evtR9AvN9d/pTgVnZzw2mWIjTIHZ/g
Te42FlfxvnVjrmuwVxUfOJNz095VLahU83EGHdnF63TQMUxeK8drIrSKeaHMD+je
j+p9S7h5UxSrx3vHv5CQVYC8xQCPTtlegxZPh/ND1fKG+tH/NROnsPkVvC2nGOoh
eXQH6OZJRHuhpsc/U9rHRJq/bosXEiyRSzXlIxZnHeBoAvFp57G2UzI6Ob7qIMRn
uyV+yhPPPiNIq0IBkh+u3+R+UYa7lbjuWC0WtUotOFPs6gdBhBsVbWZuw0DVIXdP
tfZ7hZO2/Qq6ECLo888kPL1kY0Gfu3mvarKmY8ogewlCQ5ekGqxF0iiHeEunKsOu
zycm5sfWwbnqZwKdQKKHrdCkmih25J/2OLzjqGyYBHbFeBeDI2ce7nt6skRqDupO
6Md/CCaIyx/oAF1CQ4Q0plsadRgn9L42ynrz5/sS9IEVZFWZ4jOkCXluveD+QGzi
+t9kOttjyTpp++czj7TjgV90HAM3N7AZxDjNAn+PL9Gi6GK518+fA0VFyy54d9Yy
WsbKcaWGvTt1q1o7bViO7AtNuVoaZvKi9zPD/frzpyOJl+Kn6mWedz8uyL/5qLe6
JPEvXksGYrm6aRRgjIO3u5afvxcwzfbCA0qyRaG3uBMBmTJiB3EyCPvDtkZ6+eaY
iRZOaLRaRm2ZvpV8xTZO7PAFgh1L7WzNkFk4mUqxpcAiTchZIMQV4xmebw85rTjq
GvxTmmcjqnT1ehdAG0mob0JF9omRbjnfUcy80eK9U9GitD8UP0Xm7REe/StgJTr3
UeQ2q81EC0uk3NssUPw+bl2cSjc+EHuI/ilGHJUo2Lt+JIPt4tWYz+U+LMtO7n9p
6TF8V8rlf4oA9DYx7p62N4PsglQt/vmqJIaW2mZPTlrpSyUx+0uFe19vc/X39rFp
ATw4RxJJhq2HpVOTyQs2h61QCgOaNLLLLZ7HwOxQtdhtxTqGcvNGlLU/RPB01onG
DAp61IJ7A6Z/lRTAnIEriBbClBt+r9LMn7WvZn4AF4ypeyAp269MCM/NI36e9Ryn
g4Kwrz9MXdCmr7f2MB5jMJ3wc0EnyltBNI+hndvTBLlUIKL6CunaRS1qJmDoboO6
83BpIhi0DRi87ENiOiUSaRWiUS9Y+Ist1W/YAkrvPxCNDRwtxzEbg80SIslMXLqD
PjlNk2hbkpfEqbuocI2LOS443mvzURDPNAwneVOD8k2PZf22szEDcILA3C/e8KTJ
S5ua5AIbwNxtGWPigQ42czs0pASH1BsECzh2NC0jyizty13Iq5IELYKy+mSnzXZB
s6xEJfs+/lS7BZxouPEOdrYiixJCBeh6+fCCQRwucoy8m+jVe89iG/VeuBSxPJZD
N78R/aeL2YQQTYHsTvU9qZNajSIYY1NXBmpAYuvKNC2v/cTiF4dfUkf/1t0DKBj+
MCGEJ6wRElP275+HEOozNWaBKvqh8NZa7jfoEamFh/XY//lqlGxUnCfKV+9OyeNq
w1hIDPobv/HdZWf2S/0fP741iBzEpQqkGNu1D53WpyzFLjtglOt+mfpQmUOTp4ty
hZK4+UB4a2dVL+V+Z7dV5r/eTfOJuZUWYPkfnFMQbEuU4fvaBYBqoTEGSZc1kYGA
OKEaShg1AFu0ksQwNwS7Z2e2pUVjDhD7fzlP7wSdEO6tC9XHEov2GydW8JmUa22z
QL61U/81x4PEgPCbgVJ3vD++AHH4QbGUtMfCZFSo/kS2E2tJevWbI0VCUa6+Augi
MN5T/zzSne3y8iMhruT2eTusLA9ritZWmCj509TwuqnoiumdHXipyFruNiIGSXJJ
PL0erbo+rlB/if7PSkOqnIv01uhjKZuoCeqsPbIRkJGOFjow1GnZkBFDjrFtysgZ
NG/v0UbK7wAFRG7WML0L6LFluT3yH1yMY63jKJsE9yBXEqF+zAKv8f6ycf2ujkn/
J9mGwy+dfXKZpGhFu2isSZ1/Hl12vvP6LSjr72/bVXY7trEkrd5VhEBBzg9sK/FA
7VHX5HGuiJvEdNKHXTUYiE2ZIqI+Aexbky3OkQMvIiWHbDFfDo3f6Ju8jRJqq1vG
3keJIhVTpTTYnzFGzwDSVgBC8WXbIuHcxejyzTkZn8yuV5WdUhloVSvC5wZyY3tz
R7GhjqaIadErOnwlX25w+ahtBLznaB/sikxFSN64VpK5l9Hi0eof/yf/DPHWbPi7
J5SQjwvf3RAXBLmUBp0qZ9zEEDSdbbSy3Cuwr0LjTzubC/y94Hd7t9+WuH1o0GBZ
7Wz5FC/gANOseJ2co/ahFn9krI2fTBEcCbDBQrilXbU/QDt1I13N1x7dB1u3DRgC
k0gWEEb71llU6ripZjHwdp0Au/Nd6n426wSCkH6ucBy9YVinnoYt31QCY9nt6Qms
Eov9m8tbsXkYrPPOmBOo6ESsx+Xl6Yf3crTxNFRdYOyqfn0VaoEfghZuWSbfS/1N
HB2FWnowv/EK/yMfjtudqWAj3CILgYHcNyfR+otuvRjYq78gV6y1cOw0U/Yok3Zp
bUGBB8qIqh++fRxU7/KIfHo+rPy6KvPlE8zyvZjjEHMj65N/5fEkenK9jtijET1u
uD4ECQjKCgOUBoatPH3hnM+bMyjn8jktU59OYWpdb2Yw7aQqHOyfpqJAamN3AzAY
ydP4XgHbx+N2xL3fxLzswFMIrKR94L0UQYJUDgqG28ZHuM2Nl7NLjnQXvEXx3st+
w6StAZ72KwzE+7KtqQSi73Kqes4vW03FjAJWx/vtGr4MpYe7dP0PRbuVGaVi2yOS
4EhipGASLoMByFbBp1z/9KynkxyhZ3z7HrMbTFBQ2qy5WG2OmWAthyOkPMN4mI5o
7PjPhVh1N0ERcwM1NlfG0DcD/0sUWm96loan9eQw3sQBly9/6I3jxt/LXLgrWvr2
0ScNB+0HPb1RkhuL1QPJBSLQghnQK8+AOTC7sp5ugWOpCkcX/MQ+ChQkyJcSQ4TJ
0TvKJYACZisFfSuo289ZadL9y5EVazxr9UVumsTL/P6HsvfBpUwI2v8J3cmDziHc
j9neZ+XNs1cnA6a4237u25jdheZ4SIldztst+1M+qE8I5ZxBPGu2vDmv5KM8euRB
aACu06VXgN8Tecv8puaR7f7L9Ke/liEkQ7MHVzEkv/D1/dATIGsG/NcLnIQ73fsc
JTKlXJbZNoq+HxVUfm6y79nPAAzs0HGprhgUjbJlB8J8yPtlKv/dP62dbLpNaNcN
+nkIxze0XpHerFST8zqe4YKYyQO3S2nBn75qwXBnkZ6eY+lTMVLxDjG29enQ3CvQ
+5ZLS8tsr/5d+6Y0nuxNJE57/vcjdy+ZeiKl+bsouFxZldMIaxf1XC0Vhzpnqcg2
gipBOGCgHbJyuEf2/AImc0NfXWJ23BCHfjCttpAiYCahGNgqKGZEilTT6qUSC5BK
jWG7kU5gDfOWaqcdRY8kVaeR69NPwfXiGltGd/5NsT4inwR/ZeiPK5UNE3QZ3oYS
JGhqdXTYf1+fKmF4lZmOqul3pcvJtOgClJtVPA8mVRLKKW1OS0S/pFsQ6q8GcvRq
Xx6uEJ6R4JdNbW7PAGtcbu1asw3yo6K2xyne9GWeEixXDMi+WjjezZKbs83oy8b/
xwi4VEuHAm4trq04kZMxXuquVoRYunSahB7RN2LjKTS44Le5KcIe9SmtAeUd1npj
1D/x4byoRlBoGtsO/kohj9jPKzvflWPJJC5lqU4dJvCkNGw75e+PHNr3svznBpZj
cvaPyTUIUv51L/qks7VyAKoSLvk5PBp2OxdAJ/+KLDJEm/Oigx+EG6UbP4T7W1/O
RMtzPVQo7k516VulT5HoldmcriNhlhkPWxQZFD44k9kWLPe5bIDngCRlD5MM0lw5
948evS28zwj2OYWD+1LMXHc9oRvUOpep2ejqZ+OL+HMdAonBwbRa/8TeKN2Jpt74
/KJMX4OOBC3Y0ujA4EWczdC46YuoVbZHH4rsAGo1wv6Vpi+s/zS7SoCR0gJNCiHJ
hbKMEmMhGpEUPE2CkYG0aut+in65CrmWQ1zDtoVE71Iuqg2RanOzI7d+d/iF1rAS
G6CHPpDCUNUcD2w/wzMCX57yIf6r7P/KHwiHVvzH5XdCdp1ed+VCqndZ+6jR00h/
DfcHiGMRoV0D6905Wp+7DZeUafrFyFA4WD4ombjJBMX5o9pJoBn0N/y74O1boAMf
Ns8/LUskyI66HAa3nlXYuZtwLyZxrXZswCfr4+Q8fUTvMLy3NdFa2o+PpEjSB+eQ
d0f09XAxmD+pWGCm1i02yu/2jRAS6dVwoU8Utz2kpFuXjG+CWF2ceIyn0o3jG7Y+
q/H2ZtEN+J24Iu8f5XzRJDzNIthCtoB+AO/Fho+5olTTR2r+YtJunmrrMLCusuBl
fiUuCBlmxL4NPMmDxv9dC3LT51ZvsfoBYotrXvoWBa62emwe1qt5+lmfjNNzv3EV
EjKi7VPIsGc0NdRELatxvPg/4ZpAiGwS03P+BYQ23D998VWKV3FA/HfhwItJS41C
CXyGurplace785s4aTYMok2hAm8uhG0bNpVkJbdSYNcxOCSiVmEJEkkuwOv6WL4p
jTuC7kz5h0IQzuG9qj3xwzmaLlzjKfSVLaveKzdZf5YcqSdO05A4dxeuoD7MoJPk
bmNeO7nXu59qdKb0EhtEjJHY4z/auoH6bLt3k1PVwY9x/ktW1GhQin7NEdXTmeyw
7jWQgpo42PIwnjTi1XIAACIk6OV+335jtg/ko5RIzdDUSIJU2C6sw0MFlkBwHryc
9jh6sJXF/ITWRiAJ6D1aky8X7e/Wz2ZhXCQPsSa+/E9rTiDM2hDLwiHnbhfaQQ6a
g5tsSsZNMMWKDUzoRadRZQLFDyAd8gbq3EEXJ0Y/ymeAUiv9/4t8EG/Zej5Z2hHd
cRNIuZjw4cnDYxTmjGJO0xOSaZL/Fjw/JHtzKLHCEK0b4ZznWQy/QtgsTHFaP6SW
UkOBnSGedLDe6yJSPVBnpL9PGNfdjW3TBPDVAMmdXw4BZwFE4mWv0vmyfmFp6Y7R
QGCXzwAAeoy4F6Lh+Jd1hPJM66EUCRJVhXbG0CkFRYzN54VosiZWd4MdzzSyrPQm
iH6oBlaIaAoF5DM+fC+HbkTy6hMss9Hi2eGrPHLqn4em/U/qPPBZxlPw21chlehf
9DX0w0lxG6pQcpeegUzSzgOrGBG2pt2RrvC4Xb58G+8z7KGlu+FUecjbaxJILuxo
b21mm79Sp19sIVJxPQt47v63ILHO0AYCENGSp0RlR3CK50GSGwSEM0A66PcoqUlM
o4ECrsIcJCR+DxxvEEtJ5rbLo1g4GqnehJ0PRMAdf/fAJC1tCSV0luN6yfqcA9uf
G8NnchHhgDlpS/dalU9cnJ5DcIFumjtjwOS2D7M9A7S44CzutQg0adbxtVt1EigW
ScceWvhSTHds9FASZAahJ0Y9XCNFhoxLmQ49McuvDDHBI8+56qiXAUTaZ2aPT1pa
970CRuP93X5W/9vd273glcaqOWaOaAkBvlDCYiYDSvZ6nqcBaNjU3wLiIzv7cjSa
boHEz2BN0ZVFMN4aW4iBvYiGUaVtb2yErdW5JoA3ZCcXwx4CZ84hOLTDnXnojRCs
iSfZkQDQcJuSDDk8yy5MpNFiGmwRNjPmT3jpeTQnPElKLB8wrb/R02PJ0eyEqWXs
ssok2bK5+Wbd2+lCbrRBGwzQdhMcBg+ux1PV+P3kupBg9VUq33WshgHqoQQBF9YL
mB4tjjx3rxhG9iguSsEFTK3VvSkrodPVmqWrZpsMvRLnrBOUeHKZ8YxEBQosuhbT
SLEL70v67RrY/+pOgVhn5XOz/9Ff9NyKAbuuUSGP7YTyytS9z0B+/NUhQn4IQk3s
LWG0cdMgdH6C70BnrRVAgW7E8vjvVW9NmUVKd5Qb4hFiMFbg0XRdmEVS/qfttR8f
275i1ZpPyCf5qRKZ4/CuJSxnCOzCvhu8qxNoFouA1Xa+Y2zByvfzW3MT8XpAedu2
2hNY3cfbIjo69kOe/OEqO46TkjHRz+5eBws3+n8pxjVNct88bF8hOif7UE0zEYVY
afsqNxgXh76UpG17Nw//rKoUPvRvOymOnJcIwbNnyV4K/iddODwJgotoi4MiiMwX
jQoH+NZUaQrwvL+elY5ZUSoS0U74mq/3toegguHXhLuVx1Uh1R5YZ0/rSvc+rlId
SlKAeLbqPHmIv/cfMy/NB/wBWmdfR/PlsWSrQODTc6MrD+t++/z1+TLnqyGgWgCX
3kG0I8LApFdvvncPnBtVBcAO8IB41sfheFf0ws9uhd+xZ5l9lou0hIvZq7ONQsdF
dqIOjSj7z158c0elIaNj/A7xmlmjnju1ORIVRZVsi0qnZNFdWYS4JQyYdyTuglfv
qDTwhDGUaHgrbD0yprM9zq0dP4zCNvNkOzxRV2Ua01ebobyaAzwjA80oB7q+w1M5
Rj0p5Lywhj+9Q3pw7r7eQLnncx0K/Ic7rJ1hvqJD+wligZ45umWbBqrNs6h8l7NE
SMUb2cZW/W91jAVQ8ZRL6and0JgwhIAZDBaem2irPon7ErYfVwfZq1Zh4EkEk4AH
t2tP9J2S6Vd3fQrvnrv5J0qa3EagD7PIOciqAgsQZ49vcfVViFPZA+O9wBMt9QEq
3p8fNoz0unXrKJ+EltzNmvZrccowFmKmf6fitr2cCiezoPFpd9DOiSV4alFkRBhz
YYi+82wRWp4aMJCZIDgKn6E+greV4l4kXDBsPXx9t8sbPcAxYfZEKmN6TQmjRqoK
Er0Bq6sCuu69sPZKQa9/fj89qNYnwQQplj3KCI4OlAlyVTlDaAsISaKXpAXl42cK
ytPv6fqPBKCQJCt1jiRb4RDK/rHsa+9f7Ii+jg8ujX74LkZ9Ml43nKfPiXtb6San
naD9AbQXaR/HWePiDJx3Lf5kqwAHq10TSjFzy42I9t2ij7gcOTTTDVt5H0craa54
fkmVEBiGtcfYiCHNyQ04ftW0VssqhlNrqjCEN7sxjrk7LFWbmBlOuJTEfK2XTwag
EKUPbhuzEJPKzoslxSkc8ssu2C4LjByILtS/iFygUdI7dodl4sVqjOQdo3gSQzFU
t0+89PPW1EZO1B0+HYKNm4Nv2s0mzjzEHbZnHiMv0DpHE65yJbCUrNh6a01EmZaZ
aINJVgAfrJ4xdUZ8LakMeyz5/yatxzxfMmWfRclk59+WdURpzwbiZpKG1Cw0oJt4
XCA1vC0AnNywNIPy62Du26STmpWOBrpCDLbebQDi2rlx0D5Ux3aC/WcxslWNizkB
yS6KdvRk4t3C83Pw/3o1yuOnF7tpyQWRrFe6aqpwmuN8YGH5q7TRpR5+g55VijUz
M4pEdvS7f5VT8N8V/MdLcmjhOP7HjWSjMtkSazXQaJBRLxtYK3bpAWFvi1/uLTBN
mermpN2jpVgRilsqjqCu0wmbf5TXCIU+an0zyo1+xwt/tbaCF5mpdU5ZnTy1+bzD
6MPTKCO44gSmJGidUFkXNlP/N6n/8GtLXo0Av42wd+Dh4ooaHp7klFNNmPDa3Ebg
Uq3jnJuV6xjVpPbssPlRWIrv7ZBKav0qz/wN0lRbt2GIEEo4L6Rx5VYWEXEJGMrO
9eBlmjNlU0mqRc/57SOlYB+AYpicxHpRA1uLKNtM0cHpwSDhQ2Uvhikuur5Sd8Yz
Y7JkkLNO2S3yzeEFHXuDlYQ/3g3xoiYD0bmlw7htkBy9tupkIU5jeANdQnB1LmKD
1ExY9ycAWr0liqkdBR7rbLdO8mca3niG7KyciKNokYKbqaEjB9uZuSRkTxZkekeg
zOxetxJoBaZPpxCHb3FqfqgrEjkK08RdR5Eogeh3ZySU3QFFEgW/j0FfzPlII6Qz
lmM7NT2RGXJAG6zPYEGiIopmbGronzNHwbZLgSSPyG4wBoR808LpF5Asq47zkgKB
9Sp3jQo6hDysSo+z6HwHu7o96N90mTzhz8b96lPaPCHH2+VKUJiMvr359j4hpqfI
yUmPyyqK71JGxhn9QOX40+Zc8bG7OH5x1BcAFdkBWRPm98tY3Y+zO4aqYr/ku+La
c5XZO4NkuGWFxJr8L5p+sCjhRVTnXQYCw9o9xDNeEGZTvb9t3S5gztSEk37FL9dP
b7/61FbY7Q2TVj/affrmPrwzRdDQA2GHycmhcEG4WZWXM88nzmI4B7K8cXB94Ji7
gmbnUPWuNW4C3eLKy4MF+97EDIOGwyyNVIHhAXfX/IBDBpyuUleS9VQkal3/9mOy
sT0hTICD0JKfB4hK7inbk/76Ka/Yf445swqZmxhzo+PW1B5URxAq52UOUY+tfPmo
tJGIra1qNqeM3khUdfUMRJxfL7/JalbOK7iZXMOZCPYup2MqU8R+DAfvT/D7Yklz
l5G7bqMFPPVkWL2Ms7gWNxTKD796uqvqsb7UOiephs8NQnHGubK8kZvHoIHNuHAO
Bu6dk1j7wMknY9OcBcPferUfNE8DmRkdPhnJ46pGNd5xugCE6uPrniBejHeM9RtA
y2MyAetJdw/LyKRXQp3AKa8AkFkhp26MXvEA6e+yZLTNtCh05SEw8AU9DacRnCLQ
9FxNYEGRYilAZNyeZRGjl8tujtvlpWMnr9f7waBBJKtquCgC24jcNpi8o57qjPqv
3SnXOEURVt2+tWujzbaOP44eSoG7RIpxsegDQTweb7tQ8h1WXbLAC5JEEki8exSP
N74PsLKgEGWhtAxxPqLrXyrEr+m5Sc7Ah+26CwOBhrOWh+M3xDQvQ/+r5QXZZkvx
8dXt8ueaDquhd9ZxN+ljrhxaGgSFS5NGw8lMyZC0sdWcJ+YkyJVl1LBsSJMCj5I/
dyG5l3G6W07QYndc/1YbWpm/VMzcYPTkd4/hIRfxk5ZTjKTrKLErPpdWITDzWrm9
kFDMTOM3Pntzy8aFUxltrgipVyeVf1ILLGL8AwCoJP6EcLwnAN4sFhs5J7WLg5AJ
h9sAFiZL4PHAzAvGaW9NtIZtvAJ3wDQ/MKyq2Sh3lA2YcxM/AvpJYBS9Px70tEwX
sa7WusyQj0raYHXXJfcbAlxzvwo/3/1a6Y5lp+l+tzKshJHK+t4h/VZhZ4/xalgJ
v1EgoWenGIgdhm38/IsQ8fKeKe19hY7C+MXHa1MlYCnJA8oIrVjjGLVkoR8+OhcP
p6eWceIEJz/RU8EL1pUtcrF8aweCeKEf006JB8W3EF3QexEzpH2LFxti+yyOUzvX
0FhG4yeYxCdcjvO2VHPaUCkpqqpS2MouasbnJCd+NXIn6vSJfADkv5ZlVRcCVjbz
V65sevhYwv64r4OE9mZrpKKFEgQBONhSP3kNoKw0fDe6rPJ1ibRaETL5sxIwNixA
AUW7HqbmHvgz2Jp6Srq4znRP4jG0oDwSKRmM4lgE5pOMgMkbBlwsLy9giz46Vpmw
/bTlpy89arqjmEP1xOfIiV+D4P641LwCWZzuAqrvUQINXMpSxsjZQw35Nh/JwQqf
jyFCy8SRexolwFD2HIuxrgs2gKlZFYZLFw9hKiyUIhE69v/eXeFqhoDFKo7DGKAe
BCqoymN8STPNX/CGqj4bTfOwRpcxTVtsr99Ig8tNbAX2UEOX0HxpQ9/7/gtyT944
RTYDLE1gNelmwIfCAzHH0rRkYtYg6isfXdoi4DXE516rZ7zGQU1nH6LwcJ8xGNHR
u0sgvyMGDUE0bazm4T9AgHz9UdnFA1MriQ919Hld02zMdrYvBkJak7PMjteRe+lI
bz+WFoWutlaS02OyRUsim8A7HQoOPVxL7OxzUJnai/+EkjBZyb3S0NC9OKJ3YQct
WRJTzVaQ4LA6qfZEG+VXOptChZuSjDN6G/Cr4VVxwKCqq4smS4GHOiKHtjZDIt3W
1wmsnW2qJ+f2y8snjYxSJvdPM64W2Erni9eP84dVsB+OA54pd9aWTkDfYntxocoW
fxb2yRBC53+GVIAVJY/VBtnypEzbD8x1Hart7uM+UNs/uf5m/KuKG7uoPT2SAJyn
Qf5ivVqib7tEAuGkWdglLisUnoFO5w+Nvz648/mKTNicTkYCjv+BMnq/2Kf5XKVG
BgopkGCUJf9uJaI0uBPqEyBeJooGwcy4FZIgi4u3IhSvshQJrWIUosvc5wgwaXRc
UnYBblJedxqhSkx9uw87glLShPOKsVCtvZGrhXCTcgkL2FMPmDeCtBieWHI8YmBE
sFvDaW9ZVz25nmRTOx6dV6CTRDyvbgNryxCyj3yFz6U7WlGGt21TE+qTPDAZta8R
wfNqNbwpWNaldzu86Y5UclPeaxBlAwhcTx058WTbh63FI1lEp+bP0447SxpEe2eg
Chcis6V16+tIizhA9tjgGX3ZZyzvtOxZ6TSCQ2WW2cVFphckZbS0frEFDgssiA8z
9Cn45mxvcRQkNre8myIxJR/rgXxhzi1su7Cy9BW8qTALbcCzM6uVwAOdETRoL4Gr
VtEEXrwULVaeSlI1YwdL41Qi1ByGshAt4f1SnNVUi17RsOUzXW3BG/rJOMfT8Dvk
lwtDWmqnXZXaE8+CojBC/aGpnCfTE6gJCYiMBecINOrUESIOmRxwyG6iHvQJpihN
4K9LJGD1qykhQjlRvKoLjbaw1M2W5K41t4km2FpXhrxBtjLvr198DxoNfh799yYQ
f90LeqwJz6bzyluNSnBpfpqEClv5BkoZF5JS4FxgJVqn+reipfqJZnMCqlGEdqaH
aIhVBRaOxt4qjdQd8illPtHsN6NwU6hz4+KdXD1Iy9WE2uM95FkvD02gq7eic6yV
ltHer5jds9qoH/F299tb5t7+TU4dsQbONlVpQiEIcUzyXm9I5yQaXw3UDpdEe4BP
JRfcXmt5Po5e9JfsTCMIU4FEURkSFwXYjMJC8Uu1j6vutuvkHCTP8wD7K0hfMD1r
EFx5SWI+eYhBmcGG1jKHCu16VFArR+UCxXKvwPw448kkTHmZ9BSIZbP81A6cwwM4
1I3JJPPwaqec44ghxDUCUG6tBDoofX0kCYV3RCkT4oxZ698uIVTV4QSmf8spE7BT
zCyghdSsrQ1N/NQOjOFWDtP/rR87brejXgZs7A/aS4GxAcA1xkMxsACeLSgEvCfB
9PchmpAxgmFevRyRfEKiQPjGXH+rlWDE9HMNAlgrVgkx2MjjukoGLNmk3tm/78mM
M71SVc6roitPmCnMLNWy9skUGc1VkKEsfYn7B2hvzliF2KrzewduMZwYLY3ifpw6
XQATPINdadAGZyLtwEvAXT38jHtYKK5LQ4dKk9D79jnPYbHTeShSek/suHHICgip
nUR59zZKOcjNmbJQu8f7lKFJvMi6xcMBNOnNPL9iFZOEGr7PXHe8Upuj+FZtrzvD
l5napA9U98O7OjqiTUG2cu0SIqHMzdEWn3x6WrBIGFkDN/ozAIDuXS4jiP6F3HEv
ENKWUs9mtHl2qB3Yl9uekFDbf/zCq950fWlYOJOszVDHNjsVMVeTWc2y0GHw+Aq5
LcJwlmCUKHmHn0BQhbrzqg8qdxRhwztWVm/TByWUJfbSaW6uTclu39FLEr1A/VRh
JdNDXWCWDnz0Oj/9gYVaNf7iP0On6eMsIktdkyt2FDKPq+OjK1djrYBpjuDgjcYu
IYKI93kVloZOMA89M8dHtXQFIvqCF3fsdc948GNH4adLgAEsBt/9keSr14vzt98w
o6+I5M2rQMmZBLqAVW/8X92dkx/Dwqd4ZD7dwviGVbRDB1REcZBuZliIr/PHRu7C
kxZvhFyIi9b1yV1MlIvhRYpM/an96hO3tTuOXxzirA3qZsOuGjxJsIk02ypHnqzy
M5V8H0RxFiM6ZyXS5pEFpUiiUuJYgygPMpdBL7DYYbDpfzm6aQ0pp+7wZXHCEPOk
T8FCKbhv3a+/HwbmA29VrNiCW35W8dkHfVGXQnUAiC4/dVw0/DHpFL6+oJnM57rF
zEH+xqR7qLryvy4dgL+PVvV2cmZ1lrTcBiwltC3pze3aBzPBz9Tz+taIYIOuDi/D
DKbktDTBVIPead7Ax02gVNtD/nOlvg2DMvcVMaFu4LXU1FWWkccptC3+XXT4TF1V
bUHu1OfgkJOB/BjLPo7xW9NsMM3kS9Q3yesfzw+FpAZ0J8PbiyvWiKlIXzbTHir8
O6dUyUBYj7RblG/ERijK96hB876K74jd0bjwXi8fHJhsryKRuXuz0Dqvg45gUsgO
j5zxqpRDcm3AXq4fJkzikfBojS8NW16b26bztdJpCJ40FAbBNzUc44UoNqI5RxP5
m2qt06+jTac0m7jVBhEB5ALh+XkgU6emnbeobxlJSm3GjYosuoPNhp13v3DMP08P
IR+EAtqXKhzmX+xraEQpgUy2CL8LvrwCsdRDStByzZ5gOKtSpdipMrosyheldMhY
APjlhasRfTgx7GDMs6mfTkqeCynkOOo1JxMvqXvYgc79Hb10BN8EqAHEudI1tGMo
ybYDmnfAGOa7u26y75g2LSJDsM2O4tPqD75Hkki+aXy5qALNHOkHI98zUWW+vWPM
POlhb2/UD2j+4Wk43Op7UqSBV2fsdk/LSIDof+nHTv/kCedSInH93Tr/ZK3Cydqs
EB7J9IYDj3tVHtLghotgNKgmcDrs5vrho5v0kSCv9C4k65iqkiIbiKdEKNsOzym+
uJeML5gyAZzDwZCcN7XXgRv5m0tH4gAlKzPO/WnKIITWxutb622+3v4d4tf/p6TA
lWooEWF93S7fnJTw5oPeHbz4oOIqwuaVlAEcp6pEQTUGWRMxdZY0aU0KttV5A+xQ
CsrKDV2c+DRje47cXAHxQ/eVnTxOmLjoxNqNi3NT8yFOVHY7xHfE8uS817tA606u
oo1XIzLPbec8lrNkeSUz0RUeqSnvc0TPPvOykQPhqtyP/lPrlULoKFMoZb58Jc+1
hhShxRoG9WIVDR7Rzp8iK/9fbjNXbywOqk8nfFRK3koC3qD+kRECbgvxQWadopBO
RwRWQjNp63Tx9mrRFU2V66I+HarpCpnlbTsFXiMNxzmzlD9T38yelZXgRzhthwqB
u2cBWNBOiOWgsdaXwAaYhzwj/oIOntvKYSeKYpvLdhktG4qwb6o2Ck/FYrxTHl25
fr014MSM+GwDQrSjefEeaZ+FK5lKMJZ4s1VGjRFRGycd0uJmpcdJMNCOsLD34COc
4G7+Esif7FIdMMhovWA2GthPXsC1WXI62m1vD66qPCx8cH2nKYqswVEYnM6wRPDR
Gd6b7pkwoB5DuBwWOrGWFEzZPo3/HCryuE9K154XnDwuBVNOWT7I4xt3wwXA1waG
NnIjxIOX7EuMBSgzq+7qAKO3x7W5L+e2qa9MuRvjrwimyR8m3ZolDeJfdMfK4hEz
l2GfwHWTkEUIyEyyragAdP37S6h70QlRBZ5AvpoA7Rpju03Ct/YgpKItAuhAGAAs
gEQJgRhI27RURV/wnyON406bgRT8ccF4Yba8r8UsocYoUQcSpOQ8JMQXf/cVQChk
6u5CN7Pdl8MhZ0x+3o3w+WzFsVYJ8wIN0nrUNMKY9gh1VGGeqpSH8zZnfIpzsdcU
54YulksssMbJ2wAMq69qsVQImIwrQGvXptybl5XmFw4MIqNAvlV8GeuOwrgkLlds
MIz07xZoBcFvOwHAstqBkyxjPFh+TS9Uk2nHQu00msM56uDDPiYvZpodEwMlN88w
RBHjIihXP40+q/qhaHAk4wFH0dmr6EciZp5wQt6v/E5hBSonXsxSdAXVpQWmTfgc
qdkwVYZLUWX1f1zH6bzasX7ipy1BvKShU2XsqIfnFX1deJO7E/x54vku6VDFN0dE
hhEZAjCmTig5oDAYGVHlqSeoRkfEk9fBn/aNqEhL9HINHLTVCPypTaXz6TOqDmSk
fzKzF9J0UaA1rWNnnWPH38f3VYxDdUiUHTrHVOHBCiU29i9AAzD2tUrRxK56Cp8M
r7RGY4tF7HOq3+Av4P+xDt+7kfu+A405oUadxIYnoABak4epQTInRneoUcCfJlIu
us/sZRLBm9ynLztEbphA6B9GKsgWRYP8SaKO2fjgZ+dPG3HgMK72NYeAl+g+8+UA
/CLucayN/BG0c7sd5mhtBR6mK1HqSHeAD5gmq0Ex0sQI4gZ4CEiFtYhtSyzN+5MV
8b6VMCgQmvEUMa0bnwOZ9nbRoHm95w1vVjfyTZAcJLk1OWoMzL4jMyn+8G6jQvvU
KAX1yPzQtFSt6K4R5MHbG+HoO8jSb7PUf1lcbA8jB0DtO0tnMIFK+NhqRliJtVTr
VLJF0myU5ndqzCLykq/V5MfbUhLKXZs4prsGk7jrnX/sif7d3/o6gNmbNIsmiRbo
ZgdqYl5+opdcRreZ6F1xi0/gsnAyjNoTOtBQGdrXKw0Y6t0zhdxs3Hhi+AKd6RLw
OXyTbBGRqrcUE2NxxvzD5q/dwmNrbCCgWzSqYhsUCzXKNl3yClSf06aUqTFGu6Ji
ZEv2k3cxSFYiGOzJ9xzR3Md26OOV6qzd+kI4ewEkl4vUfSjens9rm+GRZA0VRqvN
ILLlzL/CxrpZr+ohXXBGsRe3XO86ZYAXvhJMFos0466cxj6v7BotHeV2pLhxww/9
k3iI2Im1aPeuFuogtiMGfHRuVASyktZI3EmvxjPjBFP4IKBF26OjrN0VsWHS0AR+
81lKDoJhTmsJTiIqCXucjcW30vFkqHhld07c6hVflTXfPM1+aUgIBk7vzGyAmz0z
cmo70ce59m1OD9ZGWhi5Ie1E7N1j0n9qBKIneMAa2bNdZtORXS99tAOa2FSW1esb
PWYicR5ulNIo93vhMLrCSLkRLgFSWR6QeGB71z2HtDId7KttxD5X1aAE9qNwJceA
HzYJliJb8kwEYj21Yi7ax7JzKJ3jRRhcOPf77D7JMXCaCXJBJb1oqHfeuS360WVq
i4PnpBelMg5K9cmQdJ1MH47h+L7YpT3edfE4HsWcaOY/pMNn34pYhGXwf04NPceC
4hNavKQagM/cGDSO7ZRWbYbJu9XOZ1gX6Lp6pzovDdZSDOzM/8tvXJ9ABFlfbe+e
jyH0Ez3BG1YOWNIz7ihrlaqJ7RyNoc16pMF8In0JCr3nDyu2DM7Mkwt7LqTdCIyA
d2DLGMBZ5Bqq4HO1x7GLZp+YGIghm4LupYP8LOVzUDCmgVHnF7XAbBazFvGp6nJ7
tvFrnZ9ZOSMn3aPT7MZdZbVAl4euA7sy26sjLjOB/JRykE0u1ZWVDsuPsoXSKuvs
38KvIrlyS+TVRL6TyQGvu/8IaV9PsfQVTxvWanDrFtraWmFmDXMqxPXYna8p05QN
+xzc8v6VHITCZC10Xg4J5iC6tW7i4+vZcWDlA9wnmYsRLX+kIm1ueL5KRmSWNBXx
nsGyJFmJGLFfJSb/Rdy9czlZhdv8s8lpUf7N84G74VasORK8juIvZBgw5xVG9VME
m4gz6SERcpmH0O2DA+eKxgf6TVPUgXoAT2kz+QOY11VIOq80LKMwq/jx/GraQU6r
QVmyy2ddTOG1PixQ9R+cqT96oolb4KaFac4QikbjUGf9iUNwmSVjKwXylUs8G5r2
sgqIWF0GIXvch1GBoxwhmOPfbQX2/HQ+RIAj0BWfU9n39WxENdnRylLT773y0WT1
TA5r2+cFQjensvhj9Y0NTWqV4Y45IzfwqhtYuokZeK/SWdQi5LWPQ4677O7ncwvq
Qs1nfs7qRH+iNkq2oJarGkJuvpVvj1dgZ68pdnh6FREEAJGEnJjLjYB/YMtA/eSg
Ol2/1MVIyIWWkiKJRKJMY9Jr77tkF46BTvfHBOX3GaSTiYTm6hgbClR2TKlVaWuz
yRmll/qg1kh0ACWPfI+w5/6fl5Jq11CnCxbUoidrTev8mcFbYwPqbJ/S8Ov9BJG8
Yb5vx1a/Az77PclelGQW80G5baMrMwZwmOXBT9x8z0xRo1fu/3U81wnjU/Tbw+Ho
sIsye8VG8N2A+t9Cg/nHHnxY3rYkxGVT3JGCFtPCwBcNYHoKtQPQsdvLAPTYZANC
U7i2bwe/F6h0aMWilfADDRD/uFRBgKPmkNxT2y4Dhs/qF8UStbmRymOCkBfilyx0
NUgv/JWCed5TX4b2hJxUmrHsmCTOd3EcL5FnSKkJaA7p27bdE6b87Yoz472Q18aP
R0yraPzU+BTTN3WTBUaVqwAhhFA7TbezOpzR/jHVSLxu1FEJJgO7lwNYxWq/voG+
sOdv9IfZP9GreQXgW463BQnRBylSeCokFyeltDFZHurZzeXhVsGkMc7I85rpbvF+
aAZPO/ovcy74COmcpgRxbr9n/49DgIwWQG1AWnh5qA7gx4y6ugm7i295kdjeP0LI
OzbBnTs0cGADoz31E8Eu+2/U+XDriVBUG+A6HlIY8DyE+reUW1U9NcLjCP2BixPn
E5sH3qmTjA4PzWI53XFCMzXV/6u6K9VgsfzgSwMryfGmum+QUBNcZN2FOdPqWYTB
nRoGdHZQWrqLi2U6BuZrmLN0OD/fpCCqyX/FD2xyupOwzyf03FOcqp4rlxWuY6eX
6lbuJIGyFc4uO8vDfLIBmHpE0Yyd9s2RJ2xzlZvxMFEOjxMEvKhj+ilx9U+MmegV
Y8z7C9LiLwj6mi2pyQmh/sWnTCUhJlsVETb7jg59E8659AyiZerg3H19JtlX7Kfv
cKw29xfaOgsyQ00EAL9HjSVzQAPXIgjfNM6AJumKx4amLc0N8KJxzMSRusCGqemL
+txVEf/8dux7EsOHcEZ86308Eva9eSYLB8UIq7UVQhSCILDY1Ax8s7o3JcYnoACc
m7OYZ+4GE08tkPryyFUtpgECfa0iIuSxfe+bKNH0nWeBtKkfIgRUiTM+smTqD7/2
EslQdWqV0EQtV3rwPs9eFKDFld0ZGfw867UX/Jkr9o269Pm9vmCFlLSwJjIUE3Fr
KhpIjmfpPzZSf1PSdb2THesqyGGjjkzq1vPbNYz4O1g0F9FrN5HsDDc2bkzftUut
8KYsOC7Vajp5jrQVGmE4nHvzY8T51fi9ec6pThPmCmRVpCr92427x8ddXp//9asU
nV3OKbEdwriqIxDFqeLejr3/y/kKolgTT24CIkGa6+sck2E+EDM4a9IZglnhY6Si
x1vAJNzen5ie028me+EXo5znyHmt40UcTIRLt8dorZfdQEM8Nq23JRBjazvezv9v
0vb/XvLuEE8WupeNsSdbC3Ott9FQZfWUftA8rmIw3KnqiGdgLYPszkr0xS4/dCov
QYG13h2hDAn+vvHRBixgHbQHpY23BSgJ3jna5LV1/c4JZXoTHdeozP6OOtkC5UFy
VJHZ6WoSnHwBjDM8BG5MCepz8XlS21UBb9M1JX0BARCUSTmuAPX7ni1AGEt2czaw
qpYcVFkB9XiZu8gzcApxt6wFmAa/zKfXze+nVjiIGe3S2Lo/xoe2ZdofSEbgiLX/
EY/JcFBjRrI4v+mkNgDXPZXDnITTSwmvRAu32epM01X7Ngym4KwZ3iiXI4GdyMMg
02WPlC13KvC2QpcMl+Xgw+4YIW9HhC2PjxMwtKgV5gcVpvCp+owcnz2jigvtwJvn
dcrV65nakkZAw/Qjno69iDzer+3DQEXXPr3HdD/tlct9o08O3/ZcwbUYrZvamNFs
G6ZUevbTB1PPpqPkQsuplA4qzsbHL3QAhaxa28GUMGKd1jGvW1WBlxu50P71vRUc
qVLcI6jzKanx68fCrPUE5ANUqqpkZXnp5VONBaI/JYJoOvsfj84KmESjqLCrVejW
ruPclz9e1PfZZ3KlDfv1Wt5Zx4HiSVGbW+GvJv958cLKgIyPcxvucAKUUF3ZhKno
vCLC7fRM86EHr8ZGpTRoD67UK9HjCd0AT3m+wfBlMFS6GciFeqLCS+eox5DyibSX
q4ik9wBmivnuQUPxNj99m8HXPVyFFTEn5NVJz1UPKlMKkCDjvRS0jPUG3aMOctmY
SY6uEDFo9rN57bPETVt6kdFIPrq2ICNFEft/6rH4KqJuPepAqmhsZ9V3acSPCfQj
5BsIEdiXZJxgP9/B3skT5UAHhDV6GHUmpEwsUExfYO2y/zExEy74oMvGB0C1f5l2
7uwmvR4MNWpCoVqM6JPd/IHQRfTw1lPKhf79q1cjpJmvkt3l4FwbvPJrwiGNPHd/
zNltVSXplEN/FKhi45DWjm+F/GErBzdfRPw9g6xnQHjnoeTc0gWjFO7WRiCjMdrh
e9XsIolCy/ZGIaQ8mMbrui7XfIW8sRCwpqVOCUyA9uT7iPh2mccpnIzHr/MFV8IN
ljvSmr9Zh/ATcObp+kgwI7EmqIrCsvW6IJjYDVc6C60EzUS8XBUUbiLlBZoHvOPX
3OZJfbCVFnY6QpvRjP4DVHKzzlyoxvR3cSqzDez3CCM7RyMNKiIGp/4lTn22Bp/M
LAy8wTlVXAsdqGynAZYLPATF5q2w4ayX9GKcltlmQzWuoj3cYZ7gaosjhOuAC9K5
OMLNoDYX0YGs2xJbF2DpfDE+f9+t2Yf1YshQfEyhEBDL8sEtAfq9lA4lYj5W0gps
lh5UNC/2Wixrm/ZGBdCF7Er6tsPexniRjF5pH+WE+qFw7sqFyfQLoFn39565IsoY
uBbDeRK7MNYFNAQzKTfgmeWBuco07fGGCNRVMsRz0AwMT4DBoGrnDLLpYssRxIEk
Mw2M7KlSQkGL523rU1ZFhjPsyGjaWtOecy/A6qYxOogD89k8thqIzQzBaayOK8di
9ortgFjzSLDl0RyAObGwCzqqg3l34aQrIesLw+H3N4gfPoe5+/SWH5/FCW70T6Jh
wBvJMjGV+DLuObMiCWGrsCoHeVb4EuvohpDkj0Ss3ebpXMIeIOni+AZ+L8JOIXo2
ugB481nPMx7A4JOTQk10C6pkP2SasY9YVf8vQaEJaKVgvqNoKGws7Xzry6KeNgwf
HQDVyVqkrHs4aAaNVxRbnf7eYhhVor6oOfsjjPS1DIAzweWgBZNazKbFcmulJDII
FKvmHCvnIdb9cmvISyCn9bfq/xQLHB8VjenaOGH10WatjDf3ZkZyICqUJM8+n17e
YyRl80a1ZsANUWXRE5tvlekUhq7/OjlRc25qDPM+KayscpZfCtynmCj2JSpB9BD2
QewEKJzyxeLxpo0tBwJUH5MVdG7T/h8SCbJLHzGDSVTXdPdBG17BOchKSPDS1v+8
Zmx+lmT2+1u/QmfFGcK7XkDoaitoFD+HRni1Q62UTB8t8ltrQFqX0Zc5m7pJkwvQ
Ahl5WrM484fJTvOHWItBph5cdE92pyU6aLSBnY4Nl4HoutIU3dH6ezmWaq9wGI/K
Gc15xLmUPydGsyeX+DXmxvUihb0VAFyHfktEdzFsDWhAYQElcNm08b1Q+uetb2GJ
t7jMvGJJsV0YbEosD5kmEwrE3fzMGd7si9JIfi6hg9DV5BOXzhIqb/NTpPej1r3Z
HW60XegSg5vJZdI3QBaZGW+f+hPsikdqj1RbuJjuj/yR6qJVfUKqpxwbL6zqe/Sh
FST/12Y/y63dwTo3ulP21+1Ykq7vS0edtJGjtW1Z+bTFcxANoJ1D+cqJ+hHVm/rJ
93Q5Y2Tjk7FG+z4et8PpnnITOSnTTdk6c6xG4GBvFyF44+p2WexUcBOIx05GMk2y
yFFlZYReL6qa/X8vrtclZb8U5POkD3gmf9xSB77lo7ALq2LD9lRPPtH912xVRmqF
pCbVNg9TVHnzmnsEPiUE1bISTCxZZo9pvapW3x8KCKp4E2sOIomEIRki2RBEsy43
eTgYQkntqY5aYUtAkgcnPEm+vyn/Iju6w46bzf7geL6E2lG2Vws0R9jZdfJhgVxG
nmRGHzo0JMQwoZ8KHudUB+raxB8FqieVqxtMo72W5/AAOtbZ2wuUp0nWFUlbkHKo
y+M9ylPoannZ6y+8/O3JOQVSk5L95TVQ6FazHySA0JZismd/3PPShYO1COBpHnJ3
MyFWYTOM04bYUM3omMyraIwCYVi34d4BkUmK+Bay+q6stXZ3B85jjbYtHuRVOOMD
pBO5YW4uQ3dfLiALe7dE98cahr2sK4KFTLGFuHHF/6Lm564m5fqa7M9sN/NEm1eN
mjHZkiq7VUnzCo7gz5+sLF/GPEAc5MAFDPmLCzozybI+eeaGywjV9hd0a9InxzN1
wrM40SaB+y/VVNtKizDNsXL51Y4/G+P51AmSS7ctXXElpU3N8yO0EHSua+PLKy6n
WTIF91ZR5l5OVrxg0bGzuCNYmFgCekcXOswSeZC0gQ8cSNZSwU/5XzVI1NMUIH78
B46AveIkA2kmhYNJVpK8mPHlxf6xaz/JVj0ppzmjUDnVCT4nfI4xmKB3pLyeDlUv
ITn4A54THKXYnNuwKem8fQ6Ii+/YQsRcyUkw3hoqnouVxWIEACleBvUVrxp5Oo78
ZJzsUq3m/B2+D99G+sSuDe44HLeFmkAXz1BB0F/dd1R7MccvCvDsiA7L1wlm2LsK
zrbo8o45jYTK3rQyoeZli9tws9ucQy5Q9cYjHI372cFF0cDRtWRV1Ym3z+mYTEXl
Ok3vsStMxGjBJPSLktZf1gVTIhl/1Sylgdhclu4I7Zerp7tmpTFI+2q35qPwDgSf
2e7SE1p4KYPLTv7c3bAgmlp/SvvOU9ItNaJprD9CKfO7m51U+ksom65YEdubXSWc
LfX9R2UJd5TdlXDOQEKYUER0gYjhYhfNob+sd3eWsQdJgQ3VBQEFTkRLI9su8/NI
fwZHBVGkfB4JUHjwWlGVKffprwysys3ocfVAcEq1GC3PmkwG+DoQE7DYK8ag9GxN
AMJB2hprkDt946OO/7G9nSHVOgXWN+SurMGRmnfSvw+r0A7P5F1Mb8YAPu+nSzA2
aSXGVszc9i9R0PAuHurYZRc6vIyYNl9DbbrW13p5+KR5Ogx/AeKqo9jfcDVpqeDW
xogwSHVC9mSFSpv7xGIvw+RoF2xZc7z5VEXWgJ/rcZbZQX4IlhnB5YkY6U55xXOr
56tjJ7xbpIobJOHXdCtB0e8O/bVuiNPYD4O53Ccm9pafkPIuDUSBelf8khitbmpn
8cb+kQmyvQMNm3sydVCVPqKY4Y8TQoSuZz/DnrTZk/rxF+9twHpjoDKZX2U/EInE
7Owdk3OrnC4nqxGxYqhcybJi4NMw+2YMT2yOhfGsQN4YaW8wsWSuXUuOEdGUlZHe
dd4LMEoFH9qvceTi909cem33PKnVEgnmIlNRANd7pKMPHuy6TBpyQsKw+UsbmdMl
dJr2zdKu2pqn7YuEakdC4w21ifw63JJC4nsxMBlOFhMagbW/KS2l4NXRyq0QWzOe
KO8ryoA24PLMezRu0sBx7e47hqsZkEW3PNxhMD/gYhRFCV0XAUUtcI99va1fx60h
DuNSSA+NbL9TIo98l6zlZuqH/MW0kGawqPwYpgVLUOBUVWyJsa5dsdsXlaJnDwpF
Ui7ezSxuwEOjlWJFEPMZCPBRuidk+Lc5SoRXuRNe08Cz+IJijvKu8AtZvh/YPhAa
1u12e0j/vnHQP/TV24op5v5WY/kZq/6UzGu6smramr9Gh1b5SbExjkppy++mzrww
1MIn8NmrwSGpma66c8iAIPKKsidX1OM4+8Nz8DyZUxvx8svus6tkcOR+2Oq24vlz
Dwpws8zGNKUV0mu4rsEnuJHoDM9DE59vS0S/afGW7fvnDfKUsQmzHN1jucU5BBCR
zYWAqkJIaxRay1vw+wx8b3Vl2WxoCvh5iUVKieLt9FPoTb/rYoLmmZ5sh8dzWuna
r+TkLhKhqmOSEii7hcoLs9chTf6u0DLQE4xORlQHrZbJjzk2sg8c4k0GPH83BALd
89ZFkD/89Yjnt4yI7AUk5Fmo+JbY/Jrb6e+TNjjyDLXPFhxy3jpyfJv9+j1im5rn
6A+h1lEs+hfigocgybeQgqXBseUhXro5aMnnqX7533Mw1TmSU51JlqoipoVfZJ2r
BxEoU/LQdrY/MeBdci224/8SdYYhaXpk76iMH52ftR7QsiZdNCpgMyKi2mfusWyx
6+NPvmwIF09xZkZ/eV1QsgTUIlDEAabqm7kbYZ3srWseCEYYfaCBzNgc1D3Rs/O9
2PWMRI8iPKY4cWWE81VehA3LRQD9mX+tYUCOAqvQ4B+TAk07pa9wtn2azu5D1ILY
AGVgoWVxIbQfryBvhTTSYpZL3+tLMfNqb/BgeQvvH/ZckmW1zYLJJeQkNLtnftBP
tDqbt3h5UwjOgkqhBGFDrIpN+j44+VDobwKAWmY9Nlf8O+jAtSKWLsqs6BSXbWQg
F4w3wjr0EOvA1A2CieYf98oiBXPn0PNXOHuTLiZcNlSFU3dIIL3tWqgtehMO25vu
C606PmZJ74K+kLcP1C6jqqDbhPg/6TZwRU+YycgyfXp+OBnzorpZhW9DyAU5UcRW
jpMbI85rrMQy4t0HKzaFmFO7OK7N+BJrpuTy5LiLH6RZgUtlIqfkFvsbqlN62iuB
ypbGQ4EmWlGE1tujzbacJFTlij5QOijS7Tl3dVQpoJ7tsr4oWM2Bo8fwcxaZvbne
RtM8Kah6RCCY8fX6d2r4YT8u/EA5bzrPMWjKbZfb9YloWEeVchDVXkYxzs0ACJjA
ZpBPwAluv9312tTdzf/ZwrR2f4vAaORonZmiyt5FDYPUntPxS0hQ3fVaN9ZKNgEz
z3mBPSdIk2Z5eIKIvYfjhs0cZEkREvK2WPhPo2KdkKd/0qPEpovwAB8nKYWdknap
B/7k5G9ruzEtvPzkSkZSKdPM05Elq18Ift1YTwywfmRgZiGNrH0h78qSIyOHL3t2
WzniBgd/RMoZmkAG44tdyLLRT2h5VMyMtOUTDJv/KojhkvmIRkZcUaGiVZSPLOuD
/zpAv6JMSa87s5Y/Nw2NMP/U+1pSg4YDw2OuVmDsX6Un3tuTMeLROgA0kbXIVEIv
lxL7+SHfR8t5FsjpYC4wsvo8lG9WFVf0e43qzwPq3a3TSYPYcASmJR1ZqgAZZ3TB
99mNdvC0ibxZSmlQYh7AC4T4TSwYdeVKES1MuzHGEcTu24x1N73D+PsAE3bJUUR4
vz3iyZUrer73s4lvdcXktlnILWCr7KTnnntgBd+BXbgE4th7eEko0Mf5zlxXQ1aB
Eo4Xc2qDsFKYvg+QH+oUqbWNHF0zieaYKEc4dZzAvRfCodgauM5Sc0Uvqo5LIUm2
nJ9S3eg1xX6TRLk4HizA4wbrI1bor6kMREfNIXytsTR3Uaz8LOK5WHVWjhoE5R2U
t6LL43yuPzxyORIzlxKhSza4qUNambtBU7XSiKOVeV/0acPcKcA+GixVHOI19szp
XYCoJCmR3RKUlAT0En7vgG8eL+KgBuFwM6mrWHzrB9eaxf9KafI8ruBePNRQn3Fl
0q+m4sTmyMAmeGRbrP9ZCGCb/Z3hANqOaRHGezmZsWKQEhj2TMlTb89iGg9sVaEW
ELHLd8YLumWS007/Zdr2uGywUnpKuh1RwCe7A/Yo84mmMTcCM1lsSLJXzS2YcUJd
0JmDLCLsfFTQo+slHVjnMosf/p7C1wK8kHpqO1HL2Iw11yw+zCDMxWtlrpbBGhT3
wNUlxjsSuYLs9AS5JvAM57OAV04ZrczU8YfVeDFQKTHMKqLUNJV+ckMaw16v6Rdl
Jf93a9TrVro3KLZ/iuCyrisM7rgOwMzrfn8ppwhvnajlUE16V7fzp7ydr1Q+aI/h
X7XeuL9lmHJk6jPAcM7yvgpMyOpqjnE+3fNZP51FKIigTOP+XtBimL/O4YyMKtOd
lM8GSqGAIEgZ2oUHItmB5BPHxNkXI5RGCKd+IzlF5lexIzL8PI5P/tOInsWzUyJU
omu2OUEKCN1IOTc91DVxAo4CgYqCnKmRL/mtCHizne+/13jetGlasaMt9HBWkehC
idKm8UamMXA9YUHxAlCZdP8p8NQofjk+0aJoRyIF4xFKG+GP7CyYjTvs+dv4eo4c
A3y+h6/8IzF8nbSR1xaqQtRcDRjb3246IkeKcqK6mMIdpKi2cxrDdwK9K3iifqHJ
39SDFSP0RRkP5fx52XdaBGZrV72jXrFZEAW6HCbqDOtiLVf/1sXveDVxs36zSXjX
JYjrkcTv11baZYWHmVK+pCw/ibnNuL2CmqLM+PMCd+cfKWj5Y5Syzn2KSnCkYJCx
rxcViJqwGzMXCQWoMT3lEvbny1wR5kgif8rbj/bXZGmXPYixbeQC7bWid5fP+hv4
gvyPUcjdqMbn0RJ3byzpVX9mzQSF6GwDV3FUF2pkS4iiwrkXMAjRJr2PnrFMLaSY
fRy28yhRpN66O7TJ3/ZdCTgI6Sxco1Z3kxgKzIHPyZOHFN4rQLT57/lp+k/izGsM
YRBlxymPUfN/FqQLqLEf4L+fY7zgoBNglMLiyMzR0XnMrRUk1br5wKRCbiTjTVbC
95YjIyLUsUASxVS72uKOCkb3m8a2ARHzl/gt/3IzcSmb5gTBlP7SIvgP0FwL52Dh
m1M11eOBZGpnjIAE0metARjXpJbTsDfwfqrELWLsH4xvL6RyrEsX+hKCsgNYqtDe
xT10z1fK+aCBT7qOQe6SGLXmhUVE/4PFMpQbqzbK8Ye9xMyCB6uD4iqD3o6SiFrS
yjald/rARb+wwdNZdZblJ3yorDW54ycfwKKmSQWVeJU69SSO61+defX1prZri0fO
Sn/iSePn4hGWxCl3QnZY4D/YZcQXnpsjDpQfHwj+3MSrMMrX0tXl/xo5dvebNqVz
4DT1Hjtryn/+yY+hpwZ2HuXxPAyaAPDobBi7j7OhcgnwHWZ+8vgb8K0gWYHqVWEm
b4pM8p1/SzjPqgANZTm3HlevwPK+znd4fPU1N2UeKvBR9N/Z7sAEs+N+PaKzMw1f
QkoTPaHz/uxFw75Nhu/3KfSf1SfYsC4zVQdn4TDl2xopwnTfoOT06EsXk8bxMJbC
Ri8D2sL6cQ+yInCqNS3E82VWntpRdu6WzUSs9/2aIJbkIURHPA5hiNo8u+/uGnvL
iuQfof6v5gK73A5oOKIYVnQOsW3u5UV0Hej4/RQB2RlKYsUGz8f6G1lHVHQaimwW
F2MjXU3US+0/ZiMKbtdCInnLgoiv39XoqZx04GUIirSqlICxIdridG6YDmWjAcEl
gPylBdI9rQcWl2341UVqMbcAcyO6RI8nyhS9wAvD9MbNH9tjoqwrsDHpBm08qVpK
noBr/tHgijj35s6qdRalf+mqhr/mMVkXPmT+5aaO/c7B8vzXuLlXrKoKIdRZEU/M
yMRDt59GV8XOoKTCLRE7hGUZ57MGnuAyZ9810btQuaJa94TgR1Z/g2NVAY+zpXkU
i8VdgK3IkIcs99kGuq6orttvPyDrCEOFWJ/6DuZ5hPjUiPSjWGL7g7zHukWGV6p1
KxidPZQ5D9mtWwWX7w8idncBbmMneyTpF1sz2PG+rrdRdbPOB/BLct33XtxyNkds
mIL1JVLFZwej6BU3/zH7FVmhiKdqEhEaOaIRx9YiP6JJ9pIdNX6KSpVBbrsi+acK
VwawNo9BvxI0nM+C2ISf/BHfDG0ndF0yhFClYEU+LjNPNUFJYmObjkJhXo5EQcBd
4f2GvbXE0hmnlm6cPIcvE2zWC60+q2PPel7352be1r22d6jS8EVvYhIpUxrgGfYi
yP0Se3SeY/DVARwYCgwun9nrbdjkS/suQuapUdBI6ZpDguLjOcTNr93Ns3BUH+o5
szG7bFNuTjBRXW87SgvkHIB7f1RRBEXJuF5DoaQIdx7/VXy1d0vXuzkQOZHFj5Tj
XL3Kh5L5zdz3LLVOgxaAH2b02m7JdwCzLVm1Vlhoi7QDkmVUu9s3wxYJ73mzkz6M
HlbEgwDDfcQ3hMjFovwMJjkMQMAfYQZewrirqpKCNgvoioVpmEFH62geIuN6ie4w
OZAbqpcq6FXxTZ5Uvy4BATrtRuGKX+nnzxBpCdkdzAe4WjskhouglixUhv56WzWK
99ePwg7f83JA2dcoyMydJ8B6le6ogD4d9SAaMap0uoP+CgynE+n8kheCLp6+VEI2
Tw59TXGwoPpj7N7HD+/bAfHcE2yAxSOSnK27OjDmRLyZfOJR/dCu1Ks3WV7jLZex
156LWNv6zRo4nJjecEUUUT7N/jeHImPUYCFvZcviRTk4zYf5JM22ojDdh4dUIy5g
zF4XEs9SwfAui7ezOfg6op7+9FyIKSuyxxJ7qnvOcoEcqaw8+Mplr4vpsybf4guT
Ucj6e9pD5cPkT0BIzWiZNA+NUcTAgo17H1+eoUAqIgl5pfXEKuahXm7FWLoWaiQl
e7cNEaejc63mdB/lQh4FyTDB7qWt9NXobOzcBi981m/t4XodqunptjrQefB9xGxZ
SHjaGuxXms6cIvlmvTTyR2wshVXpBWtJVqeJWkLzuAsSulq71qxT4CR8HYdyvc2/
bA7lNiDp+zzHI4jbqD8eAmV/BdOzYrd1ySR2abrdWuOUscW7C3xRetbBI2bVZ3a+
N36Am5u1CkKmKrGyeAKPyHqM61j37kt8LY4fV/cw/1hZE4UcQHlB4isFZJ07VV1p
5ehvA2ZuVOHZkSjCN1haU0RiSNoWEbLWbFm8Hozf/S6y94pVnNkkYvM6ioWQK0Oo
2QQ+mkEbu0yn6Cb9DtyZbh09mBmVS5eS57huIdWQRh5kUpTpX1qzU7OgJVtCUurR
Nsln2VZuyRk17sFKTi9ThtDBP3Imzum2NehoyTtYkco35x3v2/nfXFlRReXGkbmr
9gsc4RWBqbL5/p+SRXFIn5VGV3a/fKSA3GiPa0fImNpWehL6jvIW7RWonSRINFZn
QuqaRt+yz5fQpAN7FCvfQp2pDvlUbpx+gd78WDQ/BqIYmkeyM/zhsg6bQeKA19y8
gW27gqizmu5OVsbBfKXoPJ2dlf5RuUdXRzXIp2ZzVeS9JZdggRkY+hJdW99/A3OZ
LJo1pk0vq8QwRzVKPRTf5DQhpnn9W7reweingxUwrwL+5pAkDqq+95IRy4hrkh9A
oo/Ab2X0YxN0nXQPeMsE8aB0nDJ2rtzcJHfUx8MiFvp+Wr4quUYgKRtZARvF81NR
j8+cjsAmuIw8h+f0a57XYKuVKefm3JKetrFChYGooJHfXYWEeab7VRCJ4NGd8CgB
WfYxyCLzZhRJBph+5B5e3WG+Vs4m6GlHp7DS3K3dEu5l9cPiwOPtwVCN7cSGvuic
wiasDe4ssUeyZ83Jwi+Wx45OhI048puK67mQFSSq1DbdEwAw5ljAg0lxFJbOTr37
PB9RjiskXwvKRuD+3lQy8mcHp1E2JwwK8ZzFDQiCwJBuvAtKd75wwGxOns0rum/B
6ELfYOWy2vhUi5r61I8SjWChjVidcehUIusOanTwLHNORA055vxkiUSZkkpeZ6t+
iwB646cBDjI1OTlcu3LM6udiGwTopHChJTmsmPfLtc6xXdm/kTGSD/84KIUTSES3
0/hTpbKzVNKIKqspWbO9YTw6OyvEZFL0HNC16dahS+YTXg9QlAQhy3Vv3unTTk4z
fRqED+tLsxOVg9uPD8iZzoGxpntlUIKHU1UMKmo0bshyn/0GbfuIgJmq/LF1VAsi
HdPNRcb/gzH19ICfDlpXWdHKb4fvluABd2CVaEEEsCa/Iz4BqRHGmA4Fqif5bOVy
FDcMeASCMdwcGpWMoJ60o4IwwPy8ibd+YBSHrhF+D2n2+o8xRaqcLq+tMe0qMDTP
d8KqGJqSqQ6CGqFaNGj2AlBlubJjSIIKz75sAWWBj2cyp4MrOC8LPlsstewOWOKr
nNXgX18e1GNwCwHJ8iV/TH6OkNfDvrDlnR8VQH+uUfcyKtpIbK+FZihJ3LLS0bWB
Kt93A5uMEIsuF7gpT38PD7P/LG4gBVQhEAYwPj9P1AjoajkCtcTxcNRjRueSncsN
71AdpJNgDJGEDgv3AYk2pEs+S5IYmS5wOU1IQsFjVgAPLHQrHklj9w7q/FC239HO
R8JOQbeOgEHUQjsWN5yFmhp4OrQ8khg3cNi45Vg7mlmhW/PbF86WV48T6DrqCaxS
1MB0yxCaEp6MgPX4JnnnBbj9+PnjhS+nciNvBQ0cOK2HH0Nzl1kZyJbYQ9U90rAa
ruOBKNFRb8T0qhUi2cl7q6jplbY9fVSxWvOazEGBQjIT96LrYXVCehC3KCze+OWz
UABpZ4qK2iK0mP3RapxM+rjFHW6f+S/Huz3ux5AzhQfnDOgEw4rgf448RIwyEzG2
saO7f+f0eSveUuPsWYjixpRqCffAhrmO/L3MC+MXXE58FEH0OGg61T58r0dT3arw
V6ioFUo8l54Fl97hmg0ktgUgoLRK62W+NmcaLey2jBobhFOD3/6ZmltqW2g8ViRA
UaNGfEaWyMf+92IQltVuoxJBv2Bu25GtAl+L+242fR2skj3Pmh9Gw3lz5uw5RvPy
FV8vLgVZd2WVzg7l/WsCw6/dTSv18fgCHg3hI0xT5XhIncFCI+gjigWkTDgp/b4J
5+CrPdoP5OLhCbOhd489cwwbBET1OS6qTEvdGVpNzKIHxr2rFpzQCLAKH2SZnubg
ZbxE+evZj5w/Nv0nqkVsp8MTHGEOL3a+6XnZ1s8OlFrmyzPDnoMIY+m/lflTUHdf
ngRQlSPLzB0Su1/EhwJeNlt5WTO7H4NIpcb3j5OhSTXY3yLdI1adnb79p4dRlXAv
6I9WH5XLbgkgsO7dB88ZLtDyla6BCq8YA8LXh5Zc/V4CHfAGXayySHjsffcN1t8r
m9VzDMUeTcC8HnNGjMp09SxJcDlo4jG/maIZv3HcLq3WhFIrs8Yuxu1KzKI5j6lt
pQFBesil0eJLAxuEFkKH3SfrA6oicj3FFqwxew/x1/qHhTwqSSQjhuVl1N5gfoLU
5DwfpsyNnu+8YXC1oGSXCbpEvVOygmlM67gQNFLOkIIAkZbRDSmgl0iT/lPf4Os9
5K7RsCeZcbsv8CZCf8Dn1ct0/EikM+HDmnDJSCQWH0KxJFcbc4y6b30HgtazzuHb
LDEFW/ryWSntAhXK6oV8cxSAeomDCQtfwBNAnvRnuQ7jelelyf2sIvz6TG+fSGSV
aN5y/ROo+GO2qi/b3VcCKksuQdVMwa2+0f7J+L9/PKg4aVqoheEKdHNwKCTmDcIF
Tx2kNJjf7JRpjim7ZnW9Nt2D93XI1jUs7403TTzdAuVMqRbdS1Im20KzOfLpaDpB
1Y2WFW1cfIPnDPJmAI2S1RkrIZoYqEYjbFlXS10v74cMBDcAUcrJpYOBMqIGZPIs
VtKGo4ekAILLoivkb5wwCRysg/LKD/DsUkQANwnuja4Rdcj77FCyfEC0/mtaAE8U
E8E7KDmrkEWmMNxHqFV+EnNQVdLWd6/adCbwj8GIbuMmRg2JAUFJd2pKo1JDqXnK
Xse4LLk22PE8Cgg6fwY2EBTHzKOamlfoYQkiTv4lo8bmP8vPzsIthMJfqmgmbPGw
TzMgjD1Zb8Op811CMACjV9DXaoHMfb1Avol3sgth5Yx6SRZnEVquxIUIPxOAMECa
MSYRopE1r8NpOIpYfcIehvKCqZ6w0JpxohYjYVjShq8zw1i9CsSXrBSg9dICioSH
CurQTiU5MJebpBgvcW4+hQ5Zoe7ULhxOjHY5g+NaEIns2bkMlCvRYTeloK0sMI2n
7N5PQf+hujATy2ZVp1MX5jJRMjRAy+BBMXBc8fNAIbAosQiNOkbWXGmsmdM10Vqa
PhhMnQxA0k2xvGbKnVX7VJTf9XMH+lwRE/QqJMb9SKN/4Tow2L/PmKBaIjKq01ba
6ajtZlI/SZ6Ov90nEDteFfOFL0k3iLMpkhVQ5AeiCtjfRQFM4S1EghwnE9deqgWD
qpULKHzSa+mxRjPgYtgrR6lYlSayljhcFp9Jq5Ui/z87V8U0idyLoddQ/9cMUSUN
9P3NSm3V7bzHCajkNgCIXy0zBm1HLAadCaCLAoFOJRTHoG5SAbcjHRAs5BHDO9bd
81gs6jyLcwXheU1HxsunRRfeWTtJjMCU3o6gIv9F0zI5KqclpS9N2Xldc9vn9spp
RtH4M84d1ADIlrB142zlhOwB3dMoDA0uPT606+EPrTWRjpLBmjseFGryJgsLWffO
NMuP4N2yVfxLIpKgeFz7B7szo6QIyTS7lbUzBm+8fmxKknBB/jpbjLRfve9gPAfH
w/MpfZwit4v2fkXdEk46Yn03I6R3CQJmpyti13Z2dT8/ZtPlYmag88Mra6CHfKOQ
fCAYDbiBlwXEMkRj8OzCRo6owztxhRKD6yNic0TkSj/y8GSm8wkrk+dfOhx4TaeJ
cNtTtNJGqy5EeuckeFBFRxxaGPtlXbq9YldJZfNIm8UFiOBlVK7zNvr1m+VYMN5l
liw0aHZL0BzXiUQN7gEln8HPhUXG3ByS66LocNWNDPl/TTjS3NyWdTZhSxNggLGD
Nl/AA4qFVowcMazeCWWRAfxIByRnD4iu50EFQ2BQlp9HjYJA/emFw93jM5tcB5sL
oIq6rdJvZ+7CfQEscQOJTQT6g98oCKAbCcRR/8UNnxyOSqAT3Ks7U21BkQvsfPKr
t1geyaxJnNujUxn6YH9l/ovKJ4yiossmMrstxWQfTkUlfjQKvIp+0IezxPZAhdIs
vbdy7NRMQ7wM8M3wyFacCBwOKBK/X0HaZ9Q4mGEnf21dyZU2Tk+YxxUsO69WtYWh
vVFBSR8BcfbmmgVopf3LUIciVuTdqBg9mh9fEiJeJ/Dn1J0vUNFxfKPxVNnA3FYU
tE7QpkHRVaZ/wLI2SqEoYz5+Cs1JSusWXhG8cJZOjXJ37qy+/Kwwu3uCJllMFOGV
odZfEMkj5O6j/LIOCBRXcUHY1TkK5GwceYFm9JrRvX7IzdlOVpExZtj6DjB5Ih3B
2x9bqjqH8g8YcGc1FQJD3MLgdQBe/pYVaczHVu10RIsPo1H8GmNDFc5hkLHoWyAq
iMHQreMGkDzHcPev4hJ3QclqL0DqLuKd0P1Q8k6/JP7zQ0+nOs2//tf5VCm2LxLV
+4YWAF+9YSj7/CyAgHw7ykbcUMqkKHBh1i0aF7NmZsSb0nRS3714oo6AAcEH9tGF
jLtaqvLlfGoWz1XQpMWxKf3mPj+9qoDSCdMXpg3JUpU0g2VQtcKcjWrreoPbr2aJ
f/8XwUm5iY7mlBeLZJbInprwvrDtOizAJfMZZoR7CKtFezAbWBM63Sd8AQvY44Kx
K9FK36e8KHwOOzfGUO5EbcHskDveC3A9/OeIX1sqjQK9uNpab5ehEAw8c0YqeYJ1
ujDN8rr5SzIRuQOwZbFB00CNvipyLYd/laZlflpEyQbe3MllbjrXDLW1pmq+eVCl
wKxvpY/TYZWjjyfnZVPowv1u+crm0RGoAtXrvwf9UZ9dhnA+A/CsRuID+0v7OwqQ
b4vx/rCyuZuXNoQ37cpcXkhpJmhybLsMyhQ9t/3Am62StET7lgIvaxMvaEmumGM7
hPjF8YTAuLZUtc3ckYpSISu8P9dMwimONQXrwXO01unLLy9AIEFfjaBWzFf6zNWk
Pa6g6Wkm6BMWLzAEM5Xgeb+BC21jIiHVRLQvaHEHcohW4PQNHtF51Ya266sQy5ho
0xmIPW6ZkCMEyi17f3yUB9P/g1MFeSHVdwYB3twdzEluHvpnAVGkaN52iqmrxYtu
UwuMZe46QYZ8r6+P3FGudSbnWoLAacMuydSdpJrQvuEAoZB1q0/zj1GYIakAOlFq
1GeXRX89MPRLpLqXkTmNj5NSQ+AUVb0j4fVaU5bTH5/QdE662vN8fmuG9cw/PCSb
xBwqE6W7mndNRl/sDgjUyDhG0n+sHZRP9W8rbkrm2be7NL/SkdIwId/YCMPNjwCi
dgqbcqjzyMDTNw7JxNfe05Vd/t19ODNJ58eJxAFUZBD1bz43bG5RpXBt7SEyJex9
sVEAXPuDcOgJWGH/bWT8maGy6LPQRSTyWCQIOWxYhKSrWeT5NfiKy2qy4xV4axXR
h8oaOZot9BHhJ/sY1MbOupWF/3NsOU1Abo+y0uhNyLFKVzmBqcf7afbaI6STRgQh
+zu3iTnpfwKYwXppq89e5pJeLuJdac9pS9u0CvANjOKSdTSxDTI+++4O/HuM/RCB
L+14jn3e7+uxJXcqg62zy9AvExmmNzxoX6yynrx2qAO4Me30T6abO5HoGbSSEQlp
D4ItBx/USOo1ptX699nuWCEz7eskAmYHvs6oUd9KKfMeXZHuvEFf2dyWY054qHJy
0OuFB1DhmXQwzBRt39PEMmZrPvZKiKRrDYRSJBACM8Wy40/SWFE3FIXKtHejkNjU
iR69YvNM7cl6Dsb0kMdBnd9kn9+2eXzoHvRJCm4mIRA1PZ0Rq2LKjGg0X7/FlRY6
npENIid4+5ULT1xQHXAMDreK4Vao+GJi1iUXvFoxyitISj1uYyhI3OpktY4qSx/q
ZWDJRnuivl7MzaJInmBFgzN3FhWmcpNgzWSf4GhjzTat/f4915Y0J+btlKi7U5Sq
z8+dbpOzDAooQtemBtBJ3JPwXbHKnn+GN/F5Q2EOCtkY2RDPOglc1SQuopVKYl5k
lptqKHfYem6WxPmV2ALc6qd5AN913rdVqYjxpeZIDmunUpFbrfbm+WFo+XuIDCT3
8H5b2MxaN6ZQGls1Iua+vtMmPJWwB9/f+yoNVRB5dTf/JH9seiRESfkpvLv8MJHs
7dP7C5Myn3pYhZ5evbLqOCj7cUqUMsrbJfzul1/DTigMb/o7SCI/kuQDw2gDUhqQ
oTjGySbE2rvrK+wNQos+ayqcn3IJXTMwQfDY/6kCsjE1m+BAEyHWoXPbYyJaD4w7
GJ/kz3mOOfhaDWrBHpNgL9y15E/hQK5hJj8cqXSg3CMD6P8T+wtwdkxZHm5Rd62M
/BeJtpB3HHaOKctmnxa8f9blxj71foCrjUk1MchqzMkbKyyGnuDFQw3kAp5kbac+
yCw2xmkVlHVRjl5HikXA3xWJSxWYdXYJX9vSWr8idLixbmfyQdFQyf+caAOz0Pdp
Z/V2uIClsRvV/ilmbEpEhdxaUv6/VVEdDiPYZhjYXC+pXFW0zZk2OCoaP6shBbYq
+16YrEcyvFg3xXloRojieBTm1Ss6Lshw8o3UfPfUsM4tbRGmXH7h1uaZbwmOgKyY
lWNZi+15Y92BKntwmK/5vYyyqUJ9iXpM5W8OcwbJz7Bp/yPm5ARQLlZSAxslRx3r
hhoaHwoIiEl9kWDBTvB/1KxGJVugILR8H0yxnmeiK3aab3nv5TFFsfyqDQMlcT/a
iVicK6Tdf8PcqiaSqRwHXmJWd1QNCNeBeu7mx7Z6UUaH93+fJCne41sBjjO7jyx9
zRRkCYk6RfqIJt30V2j3s4csMMnTe0Z3Cv2DJjZZVwc7e/IIybrYUXRRr24VhREr
/gJDStqAfQ6KGKIEEg7tFh6LzbvwY6NlwCSp25r1l22wRF/BlYKdQkyaRoAuZCU3
fdHBPr/pvHDxJ0UbYpeLP+GkQzrZBA6zcd+d7N7kKGt/dt1WLCA6JohGppkada3l
lupSFZLvd/tTXkzZ/mbWuimdhgVEs+Foao+3eYa9PzAnGBDsfW5dHBe36ix3E8qB
ILumo/mvGzoBOIvvdamtCirFph9dmuBfm/Ze0B50qporZ4BfSPa4pos1goAnKK+z
mSkiwLwikgkUzseHrBA+LVbdSw7/tLmDMz8J+JXqHXhFlu9dq0x2RxRuVTbY9RVh
iiYprEmVmIYp29dcOL0n6PUHLQcv8J+OvtRO14RcEr2SzzNiuSWyAUPO0cH3+hSd
52phMqqoBDvbA/FbZIRq9xVRh6Nv5SKIh4rtEZMuxZNPfkS9eXYDZAxK62tURyhQ
5a1bLpaOjRO8y006206i1BnlHAF2UNOszo+/T46y6fbXXzdEOfBwA+QiAfxJVGpP
zl6yrtXVBpDrsYOtwNL9jvgO7q92XNIvP+kvFCfz7eAqMbjnH4Jl5JiUS54ka9tR
Xo6iZKa+cZAaJJRKXXMgn3i4cb+OXYutO3Q/NYNtbiGwvK5SCHH7WyE/ZNM9MhMv
Dy7tanGwWwesiTddw5v3qaA1y4AJlec0TwP7wqJN6WsXKcgZCkfC4a6V//CsJt3Z
8jI210xBdD2Icor4FxxrsZaHxNBWKM33HVhuVRGmOo8uZaEZYzEof8ADp5l+GpXX
825lCAU949M00t6FOMYdowQmInY2jeIyorD+2H3MVUrADNkhZFvcSoIp7ltoYmw2
NVbF/t9Eyx3r/7RNUorslTVbU2UIboKGwEnNUZ+MDlcRZaAWZw1jUQFg4aG815gR
mKCQVVIS1Tw4uoCXUV7QPe/dOrAVT/v4Wly0xSyco9X+WKsniVTGrWM8xAKsU50F
2tjPf7LtUZZHGygxlH4vTRQZx/bvWlKj3XB+eCP8sQpDq4Rfw3rcPvdBDq7xv85n
spmflMdIkBkNI7gf2HMmHg/Y9ZPfPBES+LpLctFqG2skDOEb/e4LDOyyLvfMY8de
jOg7fFW7ChUjRXu2YEZBsSxjys14y5ttTuuxt+Hc4weTIO4Gai7xuym+HR5tbGet
kfIAdIikf8V9EVRIZKZQFLHs3Yd/upofFybn2mNjQvUewt7YHCVGL49qMdFUStTu
sfmV5RAfVlw37DtxFB4Qb3mi+Ii3d/9ATDgQSPa4kM/7yYoleSQyvG3lXfLcliXc
erHoA/YKaWiCJX0ySl7X6aF8hGh0pqeD/1epVzs+PqLJ7Al0m4QcLdTeg1HhGXid
uEMgVX6Qpd53XYat7omzkXRh35NRQPa4eVo1yUX+sEnhuLR5xz84h88ZuRKnOVQq
w5d84qoFjOs+uY7onzkJvQSjik7hd5KnSQxQ7vZv0/3j1MloWiarnAwgAV+4Ev/y
PXEa66MdIBfcuIj/vlpmeTIqqrTLWaqe8DZTMU+gImzNCA64p4CR3/RAY6iiQG+3
ohSHAAwUMTH79Cm83ALXDAsB8uMKVYYNvRhvM4P1QN8tc1KYRIbhTN4ioCgpEuWr
O0/v7BQlqXjN2ELQv+1mc3QhYUvtTOLPB+eWoDYTJVPzdWDusSJG/J+win9H5AVl
j4wcu2fJmYcyvEyN0poihNPaoY87FqRq6eBn0rW0BlMgJwTaWsHJPzC0rSFSaI+t
s4zXZD4xHZ32baeY7ai+ks/ilAs6gMgyvjRkQZCvyHN95X4owqAa60TTkHg2NQlv
odaOR69fT2HK2v6tbsWBKKvSlyO1LZkMmKySVfGvjeJw2xLTuQUJebOWvphcoYym
ETYmDRXnLMKSq3o9pY/UZ1KTC6QbPrjum00Vyr+rMZjJBjwSgyXLjv8cElA99akz
y5lvm4kVlB/cxu2kfZWvlh1coQXV/jiIo8dUGkEt/3RGbHK6HeEVHEniYwBc7QQp
zgPjV/kq2y51F00STPs/StYMKOE1jvCqwMKTOrdUjmZNiqavoNua+bRw719UcHtt
2vXyoG/tIuDNNBFlZYlajI8T8V/dVSBEwneljX8EiyN0QFDqbXaTrXQFlv9AAIki
bcA7itnudUydB/g810+5CsE46iGplVeky2/lOZSfPDSnfyyvWGCDeZ6bSLZDW3YX
Gu9Q7iuXLWYTYFA523/ePzsOzo9ZXX0SFIULJ816hKZxj4ScFI+Mj58IFWfU6IkJ
WOjjHCAEwqwjhvd4q4OgEtB2Bidswr6AdvkpuVUBhqzVF7mhC/nNNM+ETr9m7YkQ
1TvdzdN7pk/ipVssuvU9RdJC4IQzn1cr76yvWGH7qckEHRt4f3V6A0CMC5XUAIk+
iiyG1rROmbhWsLmWsyw3TmAKIvJr8GvCt6q9i9uXI7eLSrVwV5HnuoZAS1yjQelR
gA7pEiN3esAZz7n6bk4Q1hMzgyqu5sTkybOVZ6oLGHDqBqSSnqinX6FRYRhmw3sx
nZvG9Yx0tf00l8MP+/8Mj48l5KIlLgHR2KNWt/3xMLTM5chLgJY/BNeYeH+5zXFj
BKlYXX376gbZnwnjqbJ1yDL51WSqqo8Txk8uJ0+BUaBxV+NJe8k///kPSGPY1EGu
G1mv4wym0anYuSnN1ZMb3MiL0jlze5Ph3djAv6rpd17fwZRFpmVXIrKxv/abmWQA
e/yvjfyog1XBXlvPXbzHvVlSxKxWaIUuMJYzpa7IUr9UokI1imxGDxkhRFV39J5h
//DWgHXfiXi43Q8wZjhVF2DpQRbC2PLI6iwkj/0Pmc7WUjQHKRc038SxAOrfioXs
ZLHsEV+5+FaFXQ58ByZd4ovLstjOjnhnvWsJ8x/Nrn4BT4gp15EWkXHCBXfN12Og
FAyh86MElZA9/c6QQkpWPLcE0LP09CRRWPV3GaYWqvMuhORq6jt0Hvi0RQs0/QNg
ZRUS62OXi8eTXnqOa0K6bVfOoyE2zXlPaatKmuTYxD1HPHJrLWhNbiAGLT9Vpmu3
ClMuig+iHU+fWz8/1ePozVp3j7ooUmG9uiDUW6BtMF/qWL2z+lYG6GzKhQiGy9v3
3g+Dj0EmUiDYi1nMd8eWPDPlo7fQgOv9xOK7uSbHM5fD7c5FshZNAdGWAzkvdb19
FDAv6kERcoWFEwyxiApnwgCL2LYGF03qWsXDcSYKEw7oOd33DzT4XOzVH7DqVhqb
NZribowwKqfy2TpIUUt+NUo4X9CZpTrJn9hCeNgxv0nmC9caYgD5GpayJcKRdz7o
H6TYkPXuLp4QRpNjhaGiwD3JNcBNiw5J59XBCde9zry6IYVi/6D3aqbzlCdZTgg/
MVTe+Uiwb9QtCp7qNIzyJIh6oTqsms+QLe4M8BASlXPYCQlRykakL1IdbkcK6SOE
Np/WLgwH1/hvo9ijj8luojc1XRdM4rD+DGVnmPG7ZvTABQTSH3xw/y7IoJOQyCoP
tzr0CRTMHMtLPHT/5f8sRPGIXvjZM0B7tFcaGUYkN5inkX/jT4I/GJC0VXy7FWfU
zNmeEch43FJmGDFO9x0eJySqq4KCdR3e8+kwoY1HYhF2DL5rZPDx5jkxXOHeKzWU
r8rCd6GO7FTVmbEXIH/Y+6fVQedm5I/6vkLc5px9fTUBcSqanXlYRgXULYjSK99b
Y9N5X5Vj+LIlqzVd6702YoXukIIltKebJ8yrzF26IUMxluifMWP/EZM12GQzyLjm
J8w1fJQucdQELP81Q8X7iynjbHwIK78VMx+JYm3+7d/Om9zZ0Zdup//5qtFyw/jz
nyuuL5VofM5JizrvOuYrvd0wuk89IWy8+06+IVAs9TW++F6GGIKiNXfJhQsTnO+U
m2wD4p7YJq7COn3MkTj60wRPYoc1HhsXPa1Gtb6ybsFZG7F+GV+bKBQewJFF2HLj
yNlxIQQmUO6LY2kJKyO9WtO7w6Sddo2p4gJo47V60fMsufdCMXMPmXTdpYUrbUdv
lnmA4jDqfwLJ1ojX35kWbskta7Zbe5naMpIVwccSQvaMQLq4jREoLhqpyiLn8hYG
wgkKEs2z7w1qlr6tD78x4NcqSsD3KIrwaap2SWUKdt1uW0S7pZtf9jiaanr6VBbg
Nl1hctQS3tBdyjpUp2j4GLn66aBDmFXrHS04nkDY/vgLYUIgs2dlPlG1ecPwuxGh
1oF06VXzZOXgu0MCeNgPAwI8IvNdxvr5NXE/sYLChukXvGpZaV/hfnDhLZ7fk71y
a72t9VnV3gn6Ny8oBIRuMny3WebDbfUZN0/J0GvoQgaGrD5Y5sQvOL6Ren8Q4dk4
YAtI6L6nh5MbUxzSS00uDbtbp6slONviFQHxrh5fYpy2oDrfTiAnokvPlknF/lLY
SAY9sdP5fdXKTtj0hFzjKxWxgCjXzzb4bU4uAiQM4B9HRurlIECJbWk0JJLSRXDH
TSn0Xj06AxKalsGMwfQqbNwpEUpuc74kDnwdejJ9AZT2lqNkkqBe9gbEwGCeSj1z
S9UO8m/QtNmDBrfa7hJ+xtR4sbNWHtTP25KwpWcwiyCbFE9TDSI+huP5rrWa2EUS
jKnPCNK+Q/1cjD0crWJhslauGHiCXhtqRRtIR6VFpUZIE+B3ViVEeMtI16QeIadf
2ajgarbLTTrqMLY2TnIJzgIGepUZUL/japjk3dXLgdjPGACCnJTlwGHRqYvK8N7j
w0SyahsbfvChGQtT2C+EMvxXfrqfiuKWzS6Dxzakm4K8fffJjccEtjxtvSKY7f4X
g2yqkJPSrbkrA1RLm84fO5kn5I+O4OHl5VaRhTZVJ5uMZDA3XlldmySVAFIW3yIQ
qjK8zO0gdD2AU7Qf8BZWA7ROLP9mP6U3xY8GzurY3MwitpTtcHUimahRdRNR8qpt
GqE8y1vY2k7U43I9JeIcBH7xT5B/Y5/lQzZnOPS8TTHke7u7kqIiiBPOuN1yrcrj
q12xTufLXoF83h29qnOm0Dam7N1C9c2xHBf4TVoPC5JLTEe3Sx0WCGoY5lA8tuKx
S7md5wgyz+j8EzFpakGS0I8diHKYCWs+GGbg73U3/WMEQmhfHzReS14OBY2fDdmv
sP0jSt1qxcIOsA/IV7JMqiXh0htHcxtcszY3qoVSNhOWEdVvbK3GOUAt8AmMd3A3
/cil6v8e3yHllsKdMGiUSANmfVC5lMLvGrgZgfAhWZFntixExKiJ78U2DLJjfcmZ
BCypFfChX3t2NSl6WAYjVvRtV0HpN0Xs9XyCNXIF9p6fg+yAa0v7aiWEdP87pXV6
xqWFcjdCS04rLk56awg/rZ/6mAAfWgLtYi/SK+Bw8rUl8KqKSxSTHA2TXCpLbeqk
299w0QAjSHsbT/il0NMGSjZrTdRtC1200Vp8QoN4yaC9sArjLDBZJGIzoIfgj592
NlKeLjhR94AuHEyke9u9Mpd+r9WtTGJAg8+7JLjOktJ63q+lJ93A2IKL5I5oU+kc
v2zWlQmp6Umv4mJsT1V6pAX56Hky5GlFqSmegNB2eqs+OSM6jFH/gwDeEVneeRmZ
eA9OyHjtdcKGHWIDN7pfCPzQvVuQDlxpY/aCTRgQvCjrJdfif4vr3HwF/0grIRYe
je5/6kJZjBLabAf2FJ04t+OOuL02Kk1IyHVRcpTkPf0cqPbpyVuCYJ8zO/vI4r6r
kcRcHpQqL52HcFaSqCdhbXfyFCVVuf1jOPpVVX0QKHjXa9hF3xBpTKkQIfHfyb4a
CRgWWSYuyGRQcXN24utUCUwPAOEYOHoHmBP51idA03r/sD8fHWQUC6wzpnIOwUfh
DLPubO4wz5XkpSzKk51fOIAWMT/WREZaAqzZTHjsdpm+dhcjushnPjeFRt5F/8Qr
zwfAn7bPSvDugroDHPYz2Xue4yzuYm2+e8IxanRDRj5cmQGSY7DJmumgE8thIDzQ
oWHCYit/oUAfz8z1Zfe+gyl5ntahsPjzMPCoGU/ZgA6NI+2UmlnL8ANOqf0YdzES
w6XdP3qKAXmkr5NCRg7W2fDG/+rxuwLmONGixiwUtpmFdJZIguagqmvonWQP1r+G
5ZYcU29JXdny5l+YOYMCYyC9PGYWB2vScCU6peTfWEno/BoHc0k4VJKrl4yC1m7b
51bEMT8bXx+v9UjYqhyt6k58k2PnMuH7a1CpdN9gpuJvR1nftgCwg0KcN3VrGnhL
s5zNJHMSYLIjB1O45cs8EyRpK+O+5c9KHkdY+kkU6pT+emlNHnQ9QFLwMMslMa53
Oz0S/Rv9HIXbMdPkyIKsojZVcugwp55PqxnYK0mEPYQNEUxJHPtcXdyYhXLmuIYU
OEvtVxKLZlWK+97oARnJ21wrjWdAzKqHpxF9MblqhQ3xwwGMrIAp+GCkvVM6iqqe
rGCkThP/NwDUBFKME7ShJ9FIwb/0bJBp8XAR+Lq5OHs4uLKvcpcZyYypL6nn0dzD
wFmkmNH3b2OGdbPCQuGU/dgk85v/CXZnhjFWvLtYRAX56qa9H3QHPZkgHAxyo/nP
TJxJPPhcW0bkDDCCPSmWt3XKwPKfvEZtJNNB0j+HfofaoGhlt7cOcGyALrmW9mxt
AKRg7Qt5LwLQosysspNGWNaIH1ZiehLOGXAdSpgUV4z8nK+vlOncRx05rg+H+mvx
AyLFqKAEmSH+CK8WaKJsGn4b0cMHXO8FF4eNAXsitjAlaomvip2C5hrQjsva/I4b
1w8YDC32lXrm4xNIncARPqHqA+fpmIw1WB/i4cTXFoxs60IlZgiTSPIf5YQN60T4
fUh5qih0PzYsuS/FJKH/sP8d4iTh3VEQG/DXQR38SWU6s60bzCUvGuFNd66NgtXU
3JUA87YFeVf390JIRu5bBWnfKZe6hw0H3+oXiDYV2RNRR8nOw+IOR8fkMlAo35sK
H0QXjF72Xpo8/aCfxbB4usR60HoFVi9ke+JyFEFrqCk6F1zx0ivw6nmAnaNPPgJu
1vE0D2hqrWHWvceOYhhY76iVWFj/TH0aRJ8FJQSSWEZtaOIARyMqlGtpxaxjvx0J
UXjevDK30aBI71Gbdc9rxxr+CQ0gs/fjYuN4hfKcih2VcqsL6FnR0sk6nRJSuBQp
izmvRA73ecMazsLzpp+QLYkUgSQJW4i5oFOkCs1D2T3wA6usyok+MOXV3Qy9gH9P
VzGQyn89pivh8DugoxDVMWA6A4rqkfUxlXnznt3rZHkoo5XhLXeIhcGwSeI2cST4
uGBDHbRuYCsySWmeqCofE2Q1w1n0zBPihMQhL749zK1v+9AkEJhmNbn77niSBg1n
1NEJuzZZrQcH0sECzQFTIqJ/RE3+IdVtqt1Aq5bKDzdjD/0qA2XAaR0WQHR1nf/i
WG69G/DSX+ls5Bn1MPXCd3sbjyF8IJIxZwMu3KMv3NZk1IC6N8Zq27EqpF4SpOsn
mNsxHCRsWT9AkDd1bKLvvAEq7rEBdsExaItvxsKlCeGLhb05XUUBxbLfP5Y1c6oQ
hYX3OH6x2USX13/NWJfMWtSQNAzTdFmkySe+FNUwzc5gnoSwBDn8NwLF7xcW8924
Kxqhz1+lKGEFZqXqyYVy1gbcwe4iQd2j1LNAV+7BKyNhprUxSmt6efbX8ju4syxD
x6pxuezI/GFeJ6J8cPy8d0zyAmzKTzTR/9/uqoYz7rc7KqQ+Z4zezOSd9qYIloJf
w4DyPZxo/43OEpjTv+KFSquEmlBtJ9IPEjJTsl83/+EutQqbCinipEKO1p4yytHM
UGMnbTcF0Z9jH2mQeSwXf4zsMSYZlpE39rIGjZJTB9dAl5WuV3W37DpB4Aknpw+6
b9lqhy3gFO1W7Aud1+AVu9CyCzzZLe1lFse75+IFhQK1Oj735othktFj0NDoaI8x
twP8iHFltWlVy8IbZLGQipRWK/xdqNcoETohcz4Dvgv2Ti43kNmNlWL8NXgVT+Pg
AeDWdIABJaCw5aProNnlaVsd3MXcTfs/I15poy+yPv+eAzlLbaWNlnN1Qy3wETJo
fARvg4rtB73eU//mLM37VF3nMRi8HsStB4twtPpy9V8VoqRVbKFhsYZSfLcieMJh
x3iNAG5HF9n7kguqTNryeCljjRtk2c5cBbQl4bAcHj9zfZKDoMrN2t3+NvqHj34L
ovsRVOviGwWk/JGgSYxnvqmVxDLr0num78a52J7nsqXqQHrZhSGqYrj1KZaSCjxh
Pzcm+vtSI+EmyEQEQ3il0SbAOrnRJIOtGJlF4GlB+HkbQ5KTzped1mjLBbWkzE2p
MzwpOxau6YNX8bDZ6u3d7mfFxGlubsR8nni1dENU9T/Em1Y1TeG6LTWbz1uNAbHi
LueI9CqKNK4bXYCc+tv+RgxaWRRC7VRaY0yR7i8tC/bl2J+0Ku4+Biv+V82AUTDo
AB0f9fDm3/kYcN6Jbbp3yKKvFA7gDMAeZB1Gc3qzDW4NOezTjoKlzNzCfmbtQKkU
+CPOUWtEREws9H3fHxvlRQn3iYWPsnc+ms62E8PBww3KvMtlrCOyp4ESznevko6R
hQnWWQ0RXT9trYgz+Lr6WGMzlDapGwMbDoHjzShPsRRJoh+Df56P+pGhnrKqFmLD
c627KGpi9XGe3frGEMMtL6X3dK+OKNs02GFpCRmZs6Wf0Y0qDREsZR6UASsNTcI9
ud+bmkb5AfNlGDPSZoTE3GeNvM8d6ibYeL3rBLRQRn2FOi8ndFYTZNXYCvoMyvKz
26JUQWWLN7j67B+pEL2gxNhr2ujtvBgh9lelU2Xxho0yX2S9g5f/N90OP4EybCtU
nG53o+/HYWjdgBxtCQJvfkd/j2B3aiYtJ4+QvlVZrDJ3xdm4f4ccRJukh0Y/PMRc
tEa7bx6JfR4s5wvojb2H9rSoq9AP3AAERlj5onRC6DgbeVwmu1mDLWX/nptGIY5o
I3cM1f77w0ZhxEQrO3Ik9O9aCB5SrqhGtmlipVfzGKYtUcHTAVH6Wj55PdzYmg3Q
sPUnG1OnmB4iZQzjXyqUxRJ0XqASvxpZGty0LEESO2G2sx+TAvlNTtdsbe7oYK0A
oXvjMOCg7xB4JVhia4nPu1La7dYZTotDx/fVnK6MBhNie3YMkN8T4+D/2ySl8jAm
bHnexbMLUosdq+yeI4xRLSHRV2/mh4vMNbyZEaDsRV/dRdNoAIvkDwvtaixpjTe0
E/RI8yQG/C1i7Qyrv0Qn0AE8PFQBJBIMrvgjbKjdwd3RmVCXobifG460bV4EmG+k
XGfO/L0kULj3Kd3vDfiD7IFxbGYsr4co9HGu84q89ooUDM6YP8qIQ3wE4M+eQ976
oQs9uNiDueCQ3mvGghrnzkPw+qoWI/r4WzBhXqw0Nl3a85tvV4QL/4IYKEmyUp2c
b3QEz568J59BYhxResjcw3WvF8e8IQErrxIlZ7+J2MreaR9G09tlgAhlPsq3mW3T
hShuOgABA4HqpIbmz+UVik2cQTD/tAj0LcnE5ZJD6WMkW6wLCLxsaNhF/J15ybgK
xHR6feXMmOF63uJcub4BZ7YM4gxJKpTIeRmm+vNaa/UYeHMOQy3L61mVHzKc5lCq
4bk7EFIdVHCjlKJRBEF5tOH+YZQhS8wGhVRKRrhhM5f8QwV/HOFSBrxmdKS4hC+Q
cirp6ETPYrLrsNxXFuDJe/XE+FALaXzZI7CtkJFNcoG8Y9Icv8QmOqJVbhRkv6UY
Ahp7MfC/7na8qJVxyvqPB9X8WZ7bPtJiSYthD/MeCU1Nlm2mdI3e6Ajbdiu9s3oJ
3q74gTRmJMaZydBscEFHirDaF1TpBHVkigaGOYIpxEICQ3eL8KV0ChvGgiOaKKUK
g8G1GHd99Iyz+WAVUx7KkxNPLHz0MlHCPAAD8lB+3rWLyCznRRnOCwqKBKKdphnh
NAV8G6NztkA48l1YQcPI01BV+oU+at08llKAm//Sl5sHj7AtyDJv+TXbOLcZ4ctX
ns5GKMlVdpO/lLYXdT7IGR8J/voQvdIvesesVYZg9aCQPRwzZlLQhp2qtEe1sQk4
+e7B7b4g9hLPki+bbBehOmFwXfHMilccDKMmFqLS5Ff3ngshGPYgknu55Hlu+mmU
1qEDEaqSBs1INE8RyYdf19EvkyiIq3Y0+16zCX2vtz41Bud4Dh2T7L8M2g5ebOYt
VvqNLz0fMMYvuglXDiot2856p8xjt505JGYS4UsWpeT9pxwYyMNo9mls7y2HDNa9
9xePB1l8UYmf8p0Qy1sja6b6hcYgZ6h/Y9CbrdqMLgn4hHgtwHDQcPFjSGeXb3bl
xsSheSSFXcayNkWfLqWC3LH8Mxof+f9slmEpw1/y2EG3wt4v7jClRGfbFabJCNhd
O730AKb/x1SyDdcXByrAeeD1bt3v10oVRbaPGt2M/YL06NvKNLTx3LbWUynAk0zE
1TqQW6b9OPXQqxN32PNk7nEdxEOV4SOPvk/mFuCDDvofem6YrPt89MiFnsWoEOua
Km9wmomHCUzMmWFjFVVGRfypbagW93i/SQm+nO6wAQNzSU6grWhyDV7BRh63Uphw
0x8YmsARlErdcNvoG62/tsFeok9hXSRvJhzIEl9vcqAaawrrwW4Y7BFil2wVVdTr
l1utpUo/nddP3EKA5ynbAn8ApP0HAoo3MaoZrLrJpD8UIqMtUhfF0f9Sw2ILf9iY
bijqhrH2j1S9Tp6XnuoKA1l3Qf4/uVDPVo/+CQNbvKFNkST/Yg4P4aCRwZN/iW4Y
B7/WHGnDT3HmknWBcVOGouoxx/fBPsWaxpk1FXxALkcLS75OZX6439JkYTpYXSdI
8o0FE1UJbmBR9BfsBlfpwxn7e/onKREP5NIvAlpoF0TCbN4NJFqImpY5qWVVJqSO
krYJWzFd8DLjfpVBN2AVZ4xVH1Ac1BwkqNLlDuu4smSeSlxRtAbIaEQmjj5cpDkN
AoldCZUrBCZ+ziEm+V/e7rk4Jbx5hz0bz7vc8MKXM/XLNsbGnYGhmfTMTjio7SvL
obKpnX2T9OpD0BN1g0hhLkCFxdUGK8dJhdROh3/V1Kf80/6WnP8Xr9iZEi+xOaK9
RcMS3OsmyVqbg9pPMoGji7olOzXteupkkYfNCehXO2t9XMNCGVoQ3/dXxBVZCdCK
ECEZ4FDnhqc/u/s87dDnSP+QY4Pxq6m6XFh/p6Fku7/TlVvRsUpEZ6AHnJNp9jCr
unr+14ZfXF5Ikf5KGjRTWin2bg8qOCn1hLAsKzNzmWALKVD4bTdr6NRhsn93dNT1
r198v9/WAwsKKoq/JQa8gd1VPLZQDnZtU4m5GXFOHgkQ3t98EzCarko6muFeX3gn
jokTW3oHL8xzF4KflM+0uU/8zSlNkKt67v2EBYnxboqfXrNT8RG8T3Kaf00mt9VE
eH22stvg4HB0ddTE4+Vv7FxJhxTmcWCAOKDov5XuNyhXfVH9sdIu5a59UUTlSHMa
/I7STb6QNcEREXaBjQqOLDmLdH+kGgIqGEOdT9X4eJJ/ScI4p+5TRfYTUN3nuD8d
cGRSkNWkwbmoQkhdZamNDA6cgl2kOMdW5AD5BRn6FokgF/OIBu0UrptIdQ+ISHZD
ZeQo5XyDLgA14jN8iX8xpRBBlURUh63y2C1XGI7zguYy8kcfc+vqXg2ak+PNwOEt
eOUoC72GvszKxpK67GQVWDZk1F+QTYT5jdmMmIdX3xsDOzdS6fl8x+AcsBTq19Y1
FW1DhY72QCdUTDld+6wMPZRK2dT9pXCX1Ex8/rK0xo+6hwfsdYx3Eua3LQugj2Cr
lcKDV9YvOO2pcBMp4N+67HEx9E4ZhTAF15qwYCB6qe56GFt0XfpyXu29NKuemkit
a32IGLaiq/goAg2cay++nN6f6zGQ3IvuqsKtFa67s2/jbsyFu8EwiGz76mkjYDUN
RMfXPnaDW34Szjfv8GKSgPz93hRkMhHSJPNIuxQaR+ED7RBpZZCN109QMVxSeury
gNwS8Tayt2zyn2mI+z6e5O9AK+6OzcLriaSxcEyn7rZNEHQSy0mw8bwfH5TWes9f
K3xMa3ENHSkLGZm44F+NgxOc3vYy9xsr1/i4QtT0tfkK9M9rF8Dn2HDD4z5qIhYp
GRPNmkTRt29HDMXUhmGY7fPWr1ljIrjAGYWaEUI5dM+Uecvi/i0UvHy+aPS4I7VJ
ULnruqoA75xp9z4uUdYIlgVTU2y1jOHK3Ex0JnlNYan9AauZAVYGb1YUidAuHNIc
wCUYF6t+xCEHY+mgfKgVO3azTp6HiJgvvCgFnilDsqVV9IUJ6oWoP9WcPPvCB52u
GXHSArco6/dSFHSjsW6SFMElunZ6kFLdFqAc3FUoN+NKBAKd7RuFuc8Es3jkiQvU
icziYtmrGod1qhJCgT+eW0YulEZzYHpRXLqaJvwIxpFyjX+iZH8GO1BEiuYa+wCy
P9UgB/lGg2U2TdYh1jwUpoNs2hrdr37xQp/u4vxMiuiDIvqLWcrP5pTc2Qyh/xc4
EMi1hFeqGMtBVv9pIUtX/jZD0EOqURs7ae61u7dhzzSIQKGFQPT+d9rczqqRw0GU
uv34vYQeDjxZbedCNdg+SjYjyoC/62QK+hspNMW6MZKJZisPbXC5WW4HKk3P42zZ
PF64aBBI5qVa8On6tsHJbfhNn7kX7yEn6XMqePgK8xQYID7pRNgpiZhWFpSODupC
M7Zg6Vu+hZR6/SwuW5Bm1NCg9JngE0Waz/GHK6avCmpCGYctn4LoP50C0hXVHNf4
jt3R1qZ4G6CKXv4WzivTsmCi3e3jJ0FcWUHR7deXZRsSdZvE9aTN+8a36bOgDtgh
cGq/82AYxywncUZa5IPr2elj/QUIYyos1ppW6d9RwEry7ztA7OiVGw5tYRzLs2+m
6slFCpAHsu/6ygiB3kJuRXiWfiYpkulinKdy9p3cTOQ5ZPh0Wje4iRvEd2eNXchX
MfCPl9tZwems7cSkPiuenxHtZt6N8KorWkS4SZYQoViI0+cqol0DWUpAbiih8k1J
+vQhbQ9k7VRYx1+lUryyPO80TNplozZ+nT+oNgpXSp2EzgQJJtORwYAv1oBqkxbj
hWRiVCmUBmOZ0K+5t3GY+qC9JgzbOCZZ+XxH5IYHibYy7XrUVNeLt8CSWrZuqrzu
WYEq0H/mD33pjFvMLLIEr591zJhBBrGEyGFAf+tZZbceOZX8oERnVw5zbN4PraGy
5riyg4bBxSelJXPnDvQFm8vba65jt5M/+PC28/ulS6TpFQzlMpvDL6bZ9HPYxvpy
uanFLwpDakHa/0eYR4akI7meVYfM7MrT0sSZ5LBmBtp9YC4FjfW3QmDlm1h6so1F
LP0TBwSoPlpo/QQUfyTVPZR6FnpvZQq//WIktPz2D4v0RX1gXmPYRzJxHddkK/bO
TePFl3k+kySsdVxlrx4JuliCplLCXdP7BNBGSlXtuR5IAyBFWZsS5Pb75IpFvjHk
e4nbxEuvsQnzJMg1iMbVnC96C2pD7FP9NbD6eZuyvXfmUxu7aXpFWZP0HEKqSYbe
BZGA/jBES7QbRxzThH6qJdzCCBB7oSyhSBN9xgj3QTMYERdF8syWnsPv/vzIfqxI
IKwTKwVPI07yFMqxpQXrc03wj/PeRUh6q+rQnAWPWoZfu63qaUOKlpRD41/CpVBD
7qjJ4+LDlizFqi7BGUIbD+dJ52xOWxTJcYHFVr7qBqOVaJMIVZD9/prSMe1qsA6Y
hLhVrpJqxbE9VCON6dRaX+1XM/s/auAIXeyrudOz74XG+su+tvI6+pOJBzIODe3B
w17iSFplB4LlLZfKRthICBj/tyyrZfwAiL0X8sFLO5RFPYZktBWovfYw/iL65094
P3ed1f02H1tcLEXxAIOe1+fSA3ZH7lHXlseeOoPQB4bJs7fP/zo0L9JixVpBs3wp
vu1SuGNCNIpxKajNIneF8r30CvE8MRktZgwGaz/zRSn+xGH2t006S9CfjhvvMcYf
DLv8HO9HfN5Z62OTBSQTTQd//HKx+KeawhiT1WUmyF17+b7+82Xyg1bjoP3k1cvo
mQzdZlLCEjBbHD5egM19LvyYcxZBwVWdp5LZ2w8Jai8u4qobPdWnsWlL0QFliLCo
6odoxNUEMbriXh07u0DYnYB32V7RQ3REECIYdCU556j117aparW7v8FXI56gDHTy
z9AjXZVgZOJdJgNblbGchBbAAfIGRd+rshlaUUsgOccCzJahXGWlCfBmzkFKhIXG
bsGFvolJKkPCw3O8OWH50a/v2CjVxlDr+k5/DdzYB98HsdunBIDlm7dbAAvcQ4sm
rTxRzxTxApHEhlN6kFWEolSwOQch0zaOCSmoGhWPitX1eoFo3KgFSefU1DnR5ArM
mIQYU69RShWIK4JvQpI2aGZl9zSr81vn3Gx1rZqylsX9STyGbqNOoN7+5YoHAvzw
HJwmL7ZoWhW5yKocGmR0c+hM+hEItCE4B6k/vYOmENgRc8NKAg3sDVNY18eJsY6q
pKnyCWfK9dCY9cT8qDmlxX7NOVz9K7VO/1rQYQyXX4C4rH9203GS9b7IkPx29Zus
iPH1e/dfqqCUNFvqtrK8Db35SlLQLsacvRcOAglyzRSx9jxOEEUWMWDBvEm2crZW
+HoqZJ4kaB86AVkMGpiJfYkrAUJUkhcZXCak2qZKOGrPh0+ZoSPbU7J80FccU85S
C2vG+dKmvpd5ATMoU5twaC9RP334ed13HaPU21rZdWmfaLAVQDVYm/PNN6epK+qr
L4+58bnDMXsUZS+KVWaJy6pR7Gk7MxbEt4hu1VqWxgg04e8F50GboaQ441OX6PR1
52RPD+ZnIuzLWpHdjlLX8IMSWvkAaD3rdApAm6ie0oASOYMcE/XhSGX03yfuPWaG
qReo45Q8fTLm2j9jO9L3zIrxZ97SyU/ii8El8wm3sc3L7R9L5hJCVvfXnNKyxq7Y
2q4YKPsZrlMcQwZh5NLuv6b2TAuUBVhMtvaYbgzaXwe0PrvHIPtrPqmQ3/kOh9At
vyHIjhetUrxIVg/KRP6L8Kwa9mml3uouPTj1BvZqXXv8pgA9YBCYUXtAIZ3GRJ+r
/uaIVgS8peFwmq53K0ElENbXpDjh6hM0y8i4onpQDG4Qmk5wENuShcug5xZ9fGcx
JFt9MZmjoo6aIBDJRC/Ewjm11sJEj5q13O6ONwUo30S1FYd8CC0Y/z3Hw7rhde99
hsQws/qq1B2/ncHrB6bxH54vudQ4M1VqmWcy5xPpm9HgOmNDclfBbzAdKwcHH8uA
0pOtuciGl1KjgV5H5Q2CnlBuuAH8GNfuLEEaLrUlh2MZw7iqYShRq/TOVxE3pIhS
Z4yMdQzHaE9QV30g7i8GqO9jqyUK5h5WB3Tn2k9otteLNACGnSohbQQCS6ZnAPhT
HSre1mTZRmUlux7tRdn08R34pVI6NdFHVkzv6dzlaxrGQR4aYgGbUpwOiGNpqXvv
CKygH/IcJPo2thlJyotmyG4lUoGCxJ9MztTf7IqrJP3vsN3ZKsmD4jyTkB+75gMC
13TnPgiZFU/3e1BCv2ACIp+PAr10gJtW/2rgxvAs7dO7rSovl0W9EoyB4SfhChrl
5fyllAEp9fsKKRui3hOJ4TKfvfdEP8U7IsgYIDI5IsozS2BbdmGuKzWYuRbD9MNt
M9GJdgK3EPp31O81kXCTkixJZYKXQTaILw4gDM51PMvD3ANJPzWf+hnXPLTfa8Wc
4UBpXkIgRQycB40eQMZopGRi++5N4bEfjXgsC8lBUmzGQqRVAFopis6L47tMrTlq
Ocz8vhMyo6Xf9J5hcPABwXwQmIWz5ZEZOEMmjrO1bPUh6M9L+2iC939exwH6tt4N
EtpmrmWWcP4Cu8bd8UdoMCyna/AXxOrBZR7Ey5mCQCVNlJzNoPvo+cLeGrUSglGA
1pKX/Si3v0Cm7Lt3uArkX7hyCIv6jyk1EBOmfTFNi35M7I8x8KrUz5UExNQiFCtI
760T+QC8V4lFYC2DXhgyMkGE/s2gKxMwb7HX/5dyar7m745/l/NT9DNmtWrLMFC3
/F1EtwzlOA/ZZ2Cklw3tS4PlKPkDHCuFfirPJTJQqnqfdcSCao1zbFZNuwt6yqu2
84FPoVoTUvz7n7bZMBN7Sy8XwqWa2IHPyNKv/haODwSmCJXw/ytXMRmpBbqzKtbH
MlDDpUW/OQz4NsbID+mLLapaRVGp7XLOtnKVojPLboxTLPZlFb+V+9r3xPYnJ4q5
HU+qTnjjsuXl2xJGpLs/XLK0zxolIY6HjJEH3aRFU0P3jokAOIf9nFrIroZOrKos
mG266GAifwZYYv362p1OKxRDaGeQoynuZBqysM5+RU0Dt7LI62AqS5XHCu0rhfhJ
5Vycnfsj2LwLCR/sKCcGekjsKuELBOOBBuulD7MqfGVolKNSP1Dn+zEviTTB/aTV
UtKpehjx7ljmeMMwDRw9P6NRl2nbtv1lXhS9Ttml1tkJmWNDeiWR7Twp8HmNrBjT
lUQe5NGoC5RzQIrPDojcrorL8qy1WJOalH4I6qqxnq+8H04HlAhASMLzH25dyuoC
fpyuqeYpLVuWsMXH2+F+hao1CAvK1zgsAp3yWntdRN2X3/UgBdHDGuW8XNjOMQQE
gqklFsMhGucOBal6KyXWPBwUgLxVhl2hCSwqMaCqnphI25Isa2fjk4AG4g/pH9DO
RemfmazmLhFlzjUUSgVh4zo/PMqJretA+N+WOk5oV6GQvGgspUsYHo2bPBouvJlF
MXAinFNRZJfW0FhHXXx387sEb0nIJNFJCdSkPuOth73ylqMPYWoLYfdZvYKYtvuF
zPs56KHKKvtxK2SSusJaFS3AnxMD/KVJ3xBbON3FRv1e1k3JNoJfAxPjNoDiofYz
6sCcCfPR/1CwUPBPGQmuOrLd/dYLxjp+uuo0x8irW584XUk/5XsfGE3uBN2iKp/4
QTSYid430RNuGqfls926cxTVV4Fuip552VwbEbW63f8dazdXSOcBXc1nJocrILyO
34s4kQcDlokhb5DxZiVv126U5HysNmVkLsKasqi/IzWI/rvQ8Yd+kZqZN1X0+b7N
s4nVTEssk38yff4Yee2YMvgQmz0MkSAohSVVBQsq+o14HRyCLMZtMwPLhvpFvZzq
jxTZhbckNt+cEqLzvbohzvILL/xnYYmpH86kDX1BZY0b/YhQYT8iFDWen8TS5b0Z
R1dB5CI7qXF2yO1N/spAY9DaolTOt7R5UKP4iYVPZy2ldaS7QxJLZdf0RtrWk0ii
Q+8H1MEyIzOrQg77crjp4YB8DGniN2BMlNxeLm0r78gmfaM3ByZgWusgWLSrhqgR
3Ebz2uq7uAqubtw0GZZITQDlPR/zjXkIKaf5ZMxG3w+G8uEUqpnOdLqMtJc/M2sD
yQgPb1WaagdZR4SLqrNnslZUJb314q13JnehWbx3dTcJIPsSdwbDUH0WKlfwkQI/
8IF0Xxac1FsOWMhDbzoM99pYJVTqXxRRz0ybH2S6M72hseULf2BR1WihDPde8nMS
HMBBRKxul0MkYTe1uvEg7Lh+Rf1ffg04m6Jkubs9Fkau3Ou0wgHxuWJzAThnJX1x
/V9ScsXKX/MPkygBqGGseYrRooL2lJBOkrbIKVT8vFWfvOWMYkXOa55ubEx/LC/7
icnI9baBSd4REXf5O5s6rk7fQ/yyashDs0bFASRMli6zjGtJuav7PXY0H3RmEMhi
k11WYO9Jpy/nudO82jgiGLCOI0zgxK/ku9bogBPGTERS7Hst3Wf2bmHlTutkzN+x
XOR9NoC8ySHTts90h5hdzVm7tH7VHWwiL+JPi+wQpUxH0N6R1CmHqQZ1TaHDtDIG
WIJq/JQIPNZl4HMKRkfuKm5exLqGs2HQ9DAM3urol5ynMZYEeNvo7gNOxFikHzL5
Qcd8/Uiw3opiCljP35CgwIriYa49FB4PH9KA68iS5jt5RwGMRmLlHZO6MZLJK0PC
lIQPm2jxt2LSmbhLTh7K5gZdvOX1akbu3oUDBpWM8c4Wmt1qEr73sTctgjqev5Nb
6hByK24juYjR2HyS6MKHYRNqas2PoyTghl/rtWWK4bDKdu6s9K7zxVff3RV6oewx
JCF/mBYa2sUc5pXx5NNK7rRcDGC6MBoXdBKXNEXvDWm7i9lkG04V6ZafUIMQD8ve
4C2HQtEDkf1FpF+zus8q4SbdYdMUB+QLKkYhtMgNh5M5k6hOkqsjgSnQqLKo/zmO
C4rb442VNrbM0OmFD1v2FkEXPkpiliNpPDQWHCfG1E3dl/BlhhYAlw1UEha1m9j1
6Mj75vl+zj941a921aQc4YbGnAhtiUcAgJLV40lLEX9zqd4TBObc/iXUAaSioABl
FAJb6ZCDYNugLs6XuuJEi5jgvGMtWAliSVoFlnNPUmT0a0Sg/EJsr1vjayeR2TJt
K5aNmeBpqxFqVVstq7HxbRp9kaH5Gq2iO6zFC7vMq5GGXrXfgZMT7M9yvEVLL6a+
9p3RTjQ/5DLtskQiB+bCwZNRnR41jTvy69SkQ7ZItiCZLwfaVpvfqTgDuCPcayyT
UXVNWYm4Mf+bU49VDJs9h6NgUB/c3qIo21/mgDmQrhbT5YaIvw/PNAyBUW22PQX/
YLrqSYxmwUUUtPWBDAnGUH7wxaTudLmLyYqkgcFGYqVMoD1HarkUl7xI0QAZdU5j
6XbsDqsLCAss/rv4IjSTr8Z5mP3JVDtEDi5rmJ8cUpYI0vWywcbFZ9v6XUwWAUed
sYxo9aKRR8jQtW541oZs5DuWUqUlJL6nx20XuQ0ISbr+YIiYx7oQPDEGlcgnkfJK
shBsL4YNrze7xnCGbq4En4CGIaZ/hkKe0JbwY+hEXpLSvkXpBcaSwi+6S9p+j0X3
gZhNIWoz2+BV3L/wqq2kqS5TrOQR7UP1Y1jLzdyMwxiAnNilRhKUtu1O9PrYabNK
6Y+7wh6+PGQ5jtASA3+n/TL43vYx85dm/PwHzh80gtzAHUJ7kzyItPfty2gTAvFw
XJ9QbT2CSJ6+PR+SAA6zeO5todm8qf/dMBa+VgChcvXIjdB3n2QYVUhyemM/B+LE
hBMqi9/dPSvZWJYkaFyazizRw+Zg5IRCAPy5HkdlwJ2dmh9VDWGT1VsXYMeTntAa
4bXvQQSb/XKIl35znOttstLJe052mn0+Ngp5IOTgQzwTRxzDU+DfVSf4sGmGpTmY
buGkiOVVpKEGMK7gHijoNKTZ+ENyqMMDU7sIr5116j6WWekFuqbIByiRBEEOA1jt
eEfwfsb+3fBwXqlHI14LmXCjqFIfQpBsFAJyOvBjmQeEhahEiBh7JFvKMYBeYdm9
BSFCCsgmg8yU3ZdUxupkdoGpTNMWQ4fwFvOzy1YnxDkhPzTnc5lxAhi001i9rlDZ
qsr32lycoeiMM43Mm08SyFdRbtMuTdty/Hz4EW1yXvEHgljTv/7JagI7B1bX1AXs
eo4mQY5TZ4N/mLn2eXbmMFkktxeI7IEy0QkOvU/xK00iTyUzT2iFUtiO4Lt+Ab7V
uVi5IUVko2Phxz7qcG23SIDz77yc+YCHJNRmdsY+Ky4PrSsZ5PfWWmt2IZ9fjaeO
BnN2u+eqKlwnBxy54LEedDfWKRLV7R2CIDMEAzOuMLz6q890QhJsG6mHc1Gsn5CE
MyHPODLvD5Gnw16uRU3iL26M8c83F+5kIl3Z1rbN4KY0OIe5CcRRsXgDtx+X4EWK
w29Ux86x9026qSz2I9Ob2kl5Sr5E6hA27Ie5LYAJISwndIXNLvuc5NmgLDGln0k4
alRpWcEVot/a5XKuz4V9w0is8yWtDs9ra2pO8SrA5Ry6gITfm7+4vYwkTO45b2E7
sKDzJo/TCQ7imyZCHS5z3Ck15SVprO+XngtbJxQo665qpTYDsuUtdhkgbgDcOkac
iK7udyZp18tC7EOF6lM6ehTvE0sb45xdanuUtQNVdxK/jm3AHtT2ip9/FgHRm2pr
wecHTmU9XpgcvmT4MUGrqnYfPxyG601gtZpllr/4kR+/ZhfibA7K0EThx9TllJdI
XWFBGrhwxBUs6i90cNLRK6/Y4gDjMcEy/AhDrUfSLP1jZ+0cizH93JGUm3AatVOR
x72qHc4uC0iO2UBLzyX1SJOOt3U6YRNptm8uFKIpVnr0EBkXRxYw2yKpgRIOYmee
ALnbnwL1hTWGNiKZSbGtuVyLYSmuif7fi5lahZDjaNL9Lzznu0cIl92Lwba+caoy
g/qU4ywyM1Pj8insqTrnpn/RyNFLboELG3ikStnzzvwnqW8PNT1593Wc1wFZBEqw
08VQLb3nISVy4yE7+3dfh0Wf7IycZeZ7U45VrEelBzQyVWxOsPWaONRM4NtJ8hb2
yNCWGvJLRQZytAb5Bl+oLUzN3D7xAL40Cig6Zio7rIInRNBI0AJsc/K2RhWDX1cV
84jCX9jDJkbO/0Fi0QoBaZKzp/4knOxKkCCV+jIAJxFbQVW/fHQH80OAynPGFKNy
iOLgFm4sn42wsN4sHdcimAumOH58W2gmAq24A7nk0x+Hp5eK+vmcZlk6zXgJFcQx
Ck6ZXu6kbxTaGt8IhttQK8p06ajxyiLsAP036aQ9HgPrx7C+a9M8g2ROT5ClbXSu
h+MTOXWRBYtoKMdd2KT8RFsv1KcY6p+TyGN7JwZyuY8SvHmkz43ILnqU6x4joAPx
bVOS93oVVioRnfkIE+jEUZq5iHQifkQ/wLT/5p31IQdjjRbi2Rm2Qu7ZVzdjKrhX
5k8sfHDpsguumtjvb0qO5BwSREw/ADVSm8FGTuPL+qSwtbAmlSzHEdMvcBMNB/dV
mfXLnhnYhfyh+bhNqfuS5O8d6IBYWjJyoEnl3MwFbgCrNdFi8IetXGiF0tGoZWn5
PHmePKV/UWOsFB5orpDk1pe59NXcO5Cmbzze/QXljtYWMPbgDc/yTGodGFMWMc9W
wW8D42a3lnt07xMy/t8JbqFnQs10CforXSqPPpychuLBN0NU3F+1tzxxrYNlYPQD
KtrGtgwrDGC86IOoj/R0M/vSbt2MvQ9vDoWBqKjdAH8JlP2zJknlg2cbP28Z/rg9
Od36P4JMWZCyv0QVB6graGcsNEBqrM3aOv+IhXHq/qTGsB/mA0Sbs2Ib8+9hqFxl
tv3n/NaQR12Jwaie7z3y6EIp8jHt6H8p6Fwde6iDdwf6e0Fzxug0gAc+EaEwDurq
/SXqrUEDMfTpmgFHGdkTojtnEJZ39qDazkz6wdkRkqVlhyJ5oB69RMC5vUmZrerh
GNURnp+x1go5qP5d5Nk2tsZjWW1XY7hc6pZRuuCZhZA1gS5Qe6+fc8DRKiPHkiib
7wVo7pSB/083pq4flA6TXCtS9lTI1M5vKmshcYBMaVHUuRTKCMLWGCKRQGju44UI
RCj7GIRBOuhQmw750kx/2v3M3SF9ohpWF29Ys3rv1PJEQxZWkXIS5qX5c0DxRGea
2+kEhEUkBwPD7IWK5Gokf/ohvTO389PuvMlVcuwRm0XyTgJm7BF4g96fiJVn29ML
7NU6ygzTqsycmjfi3vTN6KP5QlKho/5LW/mcUNT/Egy1D3iaxflmbN+UCd2Ob3H8
RsmrCWPSm106/gSvVtBL/O1hev0g4zjr+xD9UbMPN/hsP0/m703Z2TmS+98iUAA5
IPHAut3uzf4cyzKencbV93r9/LwVT5j7XH8EhNPJpBGy+QzmATlmQuKzgrPQXD6Y
5cHTE6QrjwJvoWrAcEYlm2LYt0nlbNdZAE8kKbr4kMOI7/+Cglt7xaofrAgrYyVr
jkNCGtkch3dP3QjQ8gLu63DlLAKacxjXSRYniFetg8+gxKibGb9ZToAQ5pwb3SCy
SrtjfiBK+8ONnzADzK42syVUqbMQlBTQ0usU/cnwziieZYl0NtqHQPqSDLunvOX9
6TASIzfA3vzdjnBntDql20ONKSAwsQ2G/jGhsAZYveZMFEhfNQgQwL7zZqnBpbs4
JnWI7uwB20q1wqxY9iZOHRzBMuT77zZ4F5rnTSMkwHXpEZaz3aMtUrKz71q6yRaL
2D05gVXIzfFlDF/kDbwaUqfFsplFagFOJ3nPO3fnr7LQtvxVhEbFvGCaJaV0JNn+
NSjZayMA3hMA3meYsIkPMWDmEUIseodcXdEd2GD2B8BuMaDR0MXfaeDuGCiSxYwF
sLMsC+7zgw5g9Gve9b6YTIe7bqnjCBHW71STFzyW0U/+WSpL3B5dF1govo+3FUWA
fnoNsxIPxGUcAtB4oYRTTyrnIKNMtZDdtt6j0PYa/0aKdMbCD+R2LqL53do2XRKc
RJ6yl9cQQ6+q97dk4nEDE++8p9AaiW/lv777C271RmUlx/vtLMPrDcOwbgETi7aV
qMcww+kwyEcciUQBxkpF3xWfM/odnk6jjwi1RLYxHiIymXdxARUs6Lf1775eA9Vm
05j/qG5vtAYO7zZ7/xvLfl2wR6WR3Fql9+6DgOHsEAXioL1L7uF9pFH17rziWzpr
nGTgeQa6gh4kzA9qD/UimMierGQgviikFcuvgREAI6/RBeUCDQIL6ZyrgmBD1uG/
kC0BxU9NZzqXjjhcpjSPNDFFTDuwK2gbXFwVY/SOsmXvLjf0tRdovRrdWefjjeYn
Z85c0Kkkc9l0jEK5PK+gouXVxFp4ivsZiUqR7o7Z1H5ycUeGuzQqOCs3Msu2R7Dy
yE0xycgHwwmwgGXiGV3QT7JQ5B/O8b3RQJ+1oHzywc+xUOCqdN7rS5VikR4stf3S
3T/QLbrC5t/e91iRZk8UJ+lXRvbM+ycnA7xeuoi1EYlNEpI2IW6MG3VrjhxCMDJ7
TsMLdnwAR00MpNckepjwqksEIlwhf+gy1U2HSLzSdELtkpq8rEmNrgVIKL9yZZq4
5WW6ebu4UpnrNxZmSHnivvTGHbrLcK97XCi4QxagdADbrRFKg/TvwYiJIG/nEE0s
RRhw9r7ZgChgjsEHUcPDXoYyJERX9kFUxB8ofQcErqQmFWtSIxeo9XooHUrD+SWQ
H54ggxvKZ+dzJ/T0icW3mMTpfualXTD5i++HRNdgeWG0enbdhUqkag0OyGACljop
g/T6Mhr1qUSFn3mDAV0gxxKoFPNr3twgR+P2vT2X/zz66EdU0z72Bf/Tk14R2dSX
PWY5DauH2l0SAVWLJYTADnni8Gd1BD/0Foj58+7k+yC80QObzirX428yQSIzoGcS
ADaj46B9muigMsrZnca3Eta1TIgUWwglezc5crKtgzsp86oU4jtu8KdHh1eQ7MHl
zD4r0/Zy9aRM8YXF1lS4LoV7XiJ292v0hrbNTR9AX/AIvzSEkoBSwgkMbnHFOooq
yYNLXsdH+vRmv74GrcGW/JIRmFAGMRF4nkwTSU+sV7PQ4sM7d+DKGCo6CYn6IHo6
6PTh/b9fyLUFE/umzGxXRDaYkvVbfpC+HWkdu2hcW44vqjxDJ0v2Xdd1BREGUPbk
ZHZxH+Bdf7Dy9FahashXrDhur+0uV5Wq0zQpp87Cwy417ajAqBjtgx0gH5TThjLJ
xny5fypp98Qqm2ao4T0F7yXzsfy78dDaHItlPrxNTqh8e7vorj2H0Dw/E9jsKhw3
jLN8pBSYYdgEwm/c39yFHHTPYadDNYsybO0dVcWSBMkPm73uklqqfiJgHBS3AbIl
0TFBato8s57Lq4feTO9gm2DVpZwduHj667alxOCaf9S4DhlFzUqSendv1LqubsDx
WqVGbfFU+3Y9EpVOAdALdumQwgG1pLuWgJk4FEaAUBV1U8IR8xvHw7Bq7PsFoOlR
huh5rUESnWAifg4+pvDCeEi7jPU4SwOKE3UcTQIMjHPNgL4NQUPM94+MUO0gUfAR
ldxdKDLNx06IvimWmgYRoJ9efyaP1GrFJXRtaiS9N2RdJpBhFF6KTLHWwQ1KgxsK
hvoXLN7t6GVZ9KBEklY61SK+3JkyE9fkPky7q52OfSusKGo8adDTTovM1CIWGB9K
GgrXMllZyKz2RspOP4I53AwTnKoT9QWuq3g/gx5+AkQ8NsU00OGJnh0zy8TdqsRZ
w2eoSFPCx9NoYu6yrY7bIAPvxOJc0Ry4fsqwmHDPPiSoUevveBoYtfXBvepNPzpc
bI+Wlt55tdSf+b0YU880MCO3T6HvNLg/ZQ7tZv6lsA5+lR7zM4prwvflTfVEk6By
i+nEt6fr2/MNrBXG6bvCP7eXrNuIJj98knQLXbL++jU0MrLBs1UtTWMvER/edgzf
ss+6UhVNbi4ZZNVjMRi92hXniCRzdqdsFuYTtJE5jijOUHHolp9KpCg0h/EmiO8h
Myq+K0rsbc/RmAl7m51ujrgnlScm4cupzH7LFdITo7Km27JzyOQE+C9Y53qOaxP8
ruu3DmCxw8KNgh3xJ+NyLc4UCChzYZVvEKEqb+X5zh9SpNwIeD1Ks8VPv8tSem9j
ix8VwKI0zPd02on046y41fMOrH82Mba8MMVgrf8WY5XzhxuBarDM9+ZaEt9f/kyP
golcJTW/RhxYSRm6144JFADnD73aru4Jzu05ywnGvhjJH12f/oKsQkJfjlt4wto1
JcXil5rK0GvQPvKAkmfxA8FgSSFslDQ4BhauytGmIMl2C6ymqHjCAIuLqWwpse65
xPjcoFIvigS7qiZa6yBntzUuF8oRJYtDJ9NO9cfr03opFOaXTvmcQKsiO/OxB8VL
WzMP86Mcogxgg3wwnzbtYymAOrhEn1+fazsIPqBFJGM70/jxLlnQIQnCuMhpnoyp
F/N7gJIA1Gm+j2ielkMuTdjsAB84IqHhVNZCOqNsJ6IzZGpQUI+nzEmlDZ4sO/fO
UZqMFMz8H2rO91dvpD2H8HNU9txbXUqRJRQeQ1F2k2niGpHALPwB1avhtaOIGmaO
QUaUhx7rox2zTrpnys6a82uFksp/mHzlaolY8PjeuZ05oDwtg7LDaPZsjzrtdq/N
wo5gPH6FmHAlaM5ej9bkH38qX4Z44fAxamtu0tqjXpv5bUt+FZYd5o4yOVdqWffl
WPsFplYnKV5WTmcjUu2Ji2oqt7Sw67zi7kqk9zSl/VcdtTlJdPsLIrFUxuq3Qgj7
NvWxfo/cVqDYEozCpRLSliMSFY+U2jibmmSfxdlHfdFYtj0Bi8sEUtIX0Ihw/t+v
5JwGhwGFbav3gswp3g5jeu2hKt+/pk3sHLmbEJRWJEwqZImEOAOgtVl8FtpkgPnq
fJEjF4cmBD97Hs2OMqaV8sf7wJqXF0rJUJhSxLBU8jG6yqBFxrqoBkw5SeybicqA
b53aCFofeKy2zTefuzjtoVhRMWp1gx6P5k69i086PAo0b/TWpYny0dC4rQNe91Y9
QevFKRmd/S4NpfUyyQzpIp8f0PjTUhY+p0iFlVwIVw3jRVTNokCnQEGzmmtiCGX7
w5DXHxq/8v5dG31Ra3VYPoBMDTGcfjB7uB/F59FXGfGoEAm/ldubSeVzv0E7L5zc
69IkV7anMijXycTvy8m2Dr792Mo4RU5W9FNrRivjZ7a7DImbCxMNH1tA6Q9C4Rmi
D9dyll1kEXpB+33Qw2GPbMWTvcpB+NBqsFNzMv08LIvrBscp1u/ii15rbdNtfQyo
AOhjo5qbIwjYKaaE3Y48I0NVAr93/4XlCOX9dkSw5e1vFylhCSlyT7vvGt1U6Cic
DY4VdVYaVyd4/ymzyCpXoZ/NbcIepnGVHDgviLPffQB5FhtX/Oi2YBho9VzvJNbv
naSjIujbCz/jYVSqtsHn13l2B97rF4y7PbsD7jEZ8WmvUOmstncbT5g7wm3RAvGE
tAPOip5pY8cyZrhUmoo8V0dXAPJyk3fNo2v0YdVzI0UxGwaZLhDmQgR0oMw2vWdC
e4yGfeZskso5EwqzMVytrd2bdoam2p9CO6dgK6/yn6M/CCU/S+1LCMMrh2Mo9D93
wabQKRmBgEAIY1YylAeuSNlLYw1OGs3sko30RuU6M1QmMCfGBOU0mrjnFwGVX2ws
XX+Z5QQ82M0WrZXCymMoAk+I2pkAdwYWEgNc9lsILbp5pzt/Z7dEAQBzewIdOyh2
bfN2NIcomkyGgBsWPw33pHx0YlLNTnU0sdGbkJBM9DZvt37S3TJa3k3sLMx4wYCm
8XJ/XBat6WLn6fw+iLkcU5Z4dNvD3ApGUnNOs3A0cAliLlXEitC7kcb/x+g8PdEr
4XjsV38QgvjPZNtd9XcDFkCXZod1to7q3urrohJfMdvPeC7Sa/U14F38yoWHciVi
JHqY89Z7eNdaTQyXIKG/Mbbes7esmh48pvc+wEV+dmG7Q1OwxOIgymxhd9rqCOQ6
npn0mWQG8pwolVF6hVy01dRREm9JxYzK2FFXDsS2fPkGIZmebaBmlIE8SP2BYx01
qZ6bGRF26NQMtPPBkIzDli5qUtE0/0XQjddG92f/9NMyLND0CnEoNTEmzWlvR0G7
2Sip5IOFd7bi2DxrGR9vsuuJxY970vfxM3pHiuxKVM1YnZQHFgaX8dCZUPohdR4R
G48+aXf3KFgR8mZ1S4GhBsdJ1Jlt3LgLHZ6+GAKnc+V1TH635KxFGMsl8EtVTDum
oRJUfvjzIZDzCC+VIsqJcVWcfRGqSS9W7kiQ12Ip7uFg8riYB5yMiVnVZ3QtN6em
Uq0YIoFcnXILyIsA/YPHk8AlRLUUARkD+Z9fmf7RMNsNOEPk05Z2XEQpN43lUOJ2
3Ht364slSDpDLkM2RxGQtv1MtuvmNMmUwSsMVF+//sUxxZBdX1Zj6w8OCDRGVrJ4
AN62w4CW1fj3Sj5X5XBJUzA8/EUOvY5Jr3Ri1EWjAcNPABZp9REnHI9qz+scepdy
FBGe7xe2iDNWsnvJkjapnlkwi//ZOWW9pbjlhFgS6v4ZNmfyvcrrJ5l4WKEBXjsQ
Ll4OhZL+QboJ/YpCRfHs7WLDpj/DgC5qE2Jm0QM+uX4xByNk2qRUJWx7NdRbYz5V
N9kicKVN4WjSl8ijmOOiF7T4C4R5I+zMWYMhKDgP7NKQ8s8DyDTD14LMFIQLw/Iv
P1FcNw0vmAbKA5gTvuY9TvVmZ5BQu/L5m4IBzu4pqrEih79SNn/PKtfwoFlYWSAa
RkyLG+MoY6abwvP9LPzGtoYS/NdMdaNwa7/qtLfsFu8bMz0dMUMZSEEHvgaOun9W
FsqLXY5/2JRXvI7HOeNtwN6Y23iooo83FZ4vlqC3CS/AQblrwgsPC/OH1Cb4Q7W3
V86EmLpj/185TqbNjiiMcWGgKzFgMZg1bfFWCAsVnLoBwjPXx8AKtZrUEj1isB6i
e6L75KPRoed9xv6p5/xX6/YwzUkuXiUFBv4iMJUSBnnSKSeRv1fcjFfHdUbXjdE0
rxzpQ4fhOIgYnnQy+VWJ9Wblg9EtTdWrUSewaWjW+1UMJbUq3W/FWCupyuD+nTWX
R+wdrii9bU0PowKoZ4juXLyMFMxx2JBou1MOxNlqBktyNMjODbaIvpMNlR+5sUDu
Oo1VaueZRvTqfZhO8N7vmaSg33+uSUxa0L/tzgLERK7fU7Tnf3ZqmX/45uUewiln
9yEmnI4OlQD7GvUtBCPhXhTVu7bSdLIrNVrcup8qExQzAur/DgGCfYuPEjVwbWVW
lFUwt+wtCxkT+K4Z4C32Hxj3GB1TFnvmWp+RINph/gqJPF67qdV4IG7W+Y76Ef1f
reIYeSarzmO6xjlkJ/qALHFwdlgrfd8iOtUlSv/cLkSqOiCaje+NdYcbwNjdC7jC
CB8jrDXeDoAOpHrsJXAhcWKAlNzFw9QJFG/TJMKIcyz0w4G4ml6PONm/X1CY29Y7
D1M+9TwkWBKF3lhduS2ud5NRs7/seGn26dL/3PWdidh7ZvsQu3hIQRltnBtwla+2
Wb2FDspeakSS4lOlyVZEwFBiVaO5b65OtlVHZOxLerSxuiHHCA3QwMV9+nKoYKYg
GA7l2QtTZeHwkbHPv1PIfFnRz9oP07JJgYNOeTXxbqcLrOGWdS2FeFs3ZGV9xo6/
WKYFBsL3pE0OsxEyVJzk9AH0v6CydldcSNb6RSi9sYvAJs8jSEa2HTkeNUM8r8jk
gbsoPPm/pKesxCBsl/5qhOzDqQNSUlzgmLKK0oVsYRjgGOiOi21PUk6gGx7lOnqU
xqKmKazkBEMDaPQN4lxfWSXKnfxAM7551EyLhxhDcz+/YnUeo7itpY77+aQE/8q5
4GvK0ZHv0ChRGKxB0EPtUJ3BW4KsVIwJtV7sYBS29vVDAsi7oQUHxlTvaJLoE1sd
n1hqVbYedkdqlgenzkkiKwl49nySd49n1WPwhlI2bLJ+zHuBwcbD9+Jr+03A+K+n
/F64fK048E91bsdLAVakovaeCqQdfVg9IVsVu4me2l7MP/V2PVY1Ts/p2rxhz1wi
hXigiPDf9y7j7iVzYzeSjHTs3j/sALbGH7r+wbj/0E5reriPYTy1fcy/Ybzo8Rfp
zsBCt7yhiKXOFBccOY6OWOC6X6N5D9yQZb2rDeaKg7SC6db/cH3kHbhitYSLvUcN
5HXe1YQQITEoP0FcszLFBpQ6csc/+6EAvbiyvb9GbPIr/8skNQmQ2sW7fxv5fe0+
5iDh5R/bEVgCbGCb+CSkE5DmNfDGBHuvG93p9DFjFoXwNaLZV/tUdB4iNZE1lE11
EYOsJMVQAqeURL1MHslEkJHjvcoOvPYiJ2GneVhnn94yGQFkEJdBW7TRt9Tlbjv0
dHq/Zw+27kLJTus7b/UHOQvCFf0Ci1l9FwQi2DMK4no80kLpUFDYKYE4VzUc1Vc2
6JfJ/5coV5OAaR71hrNIdO/MgHPSAEjo9MAVLcJzziolT/eBvotW0UXVLcCFDAc+
yw+cNIO6tmcRnkUdQQoy7QfK2EHp0Y9T8h0WzHwqYekknkxHtHJ6tAze2P0FP2DF
vpHBbLmlcCbyCMevg8nRTJzJw660qYGBL2XggEVjW9GbEkVN0iXMWBIpliplwjqt
Dr0LIbXyRQizQIKOg/FkiBazVjfOy6DEpYACQMmtXdbhDjYf1xxKgFI/tUfEdCBE
uXgvoIY2Jy7Geq4aQHn+AybsjI5FwX8LMokVMfnFGe8fn1p7XtOOI8LBM2+NLxK2
oert386IcglzBT8IZS6Q9zthJxfDp2Eb7f6FC801r/0rwDBZK9soL0eotn3IfAO2
5FjZ3ro4bxXZmV0pZMlMyCmvtKFgLhV+TJdgQ+cKk0m841t1u4kzbSY15zH9/f1P
4eQqYb7ujKfx/AkoHFisjV2NsUY4c6duhOD9PXasnwSuvk8ZKVmEjumjIV/0jK7i
SesoARCz/Gy39d1jPyyDbLP1dthFz4xl43GhSj9qdn8dtJVQf42KTwps+0D4KNWH
wKbjrlOKl1vPow0p0aV4TzObIgPyu2vVKt188gIc/2LPCz14rvhft57kPF6ZgBid
NctVtBP3mOgck6ea3ECTNn/xSM4tjFvzLfBS2OvUcLVj2MeKl7qbxfIeVsehlogq
PXr22l31zHJ6dmr9iSvgZRQXIVqXdTh6JvoHlaGVtajlAQ1hn6hxSsK0t5flTvy+
CmKTvW4SzyrDKLanG0HcG1jNDcc0DzNpDgbTdLhqMQ6vNRLP3+CKnd8xlfOAzC+I
ynnSBcfTnybl5VMLB3LFckTnPks0VjA9BBllsjtvN5iin25I5FjPyko7+LxUY3/m
u/LA88omc7GYAJ2TyYewRUZq3MZ1DA9BL8zf7cjJMgJyuLpRqebHpEBXuYmD1iWJ
Kk80LwCN6lY+G8tVmYUgzlP7CEKVg89t+Q9nQgmXa0u+1nbC3PIE7lj2pmRIgGmr
2I4Kgd/LV1uSA/uGJYH1neZk8WAWsYT80/+NPICOv1KGSDGVC4yK3fN8OVKnj4Dl
72H5jLJ8E+Vo5/6o9TAAkWEHIFvUwib/OB6d44BthjbWD6ZNlbUxntH3aKizGPQf
tJKQwJPLln7IrksJXNkjMumDVuafIfERizgNHLJ0c8aT/LC48qi7X1DBkh87QGPY
rkBXlVbWGbtz2Xk5F59FfCj0SQPRKpSpqxn9FcRsCWHKtmBJuFiexweodDEimNDO
my3qROekO+zXj36v6tZybVXULbBT3Lb0yzS+D0NkwVZ6cQNN67jxv38DL9WGR+1l
6I2kOds4Ye3XOlgXlKzggA2G0+IDXJqBLgeef7JsP4OWiGcfJKKuI4DZtxmUn7bq
I8cioU9LKH1qLUF55ZOhrLS937FoG3xaeW0Wkw5WDee4f4vwBjzg97nhlBaYBBfz
9eAGlXejXeyQGdIHZpGJ9h/YA5TZYKKUmarm5XleMQ4Zi4lbI351ytvd1XJvJe3k
SJ7IxXXd5G/qAfphpDMjFNM7ZOY+TFue39iqjjmB/6Uuh8c3eu0E4OMWji/3rQsx
gHkhouASf9jH7Av54dBEusfPX0A6yQJDOVsXV42JJCCufUuBs0vMWsNLPl34jYXM
GJeVT3PHy1TyH4RW13bBfy7dTO6SoVheBaDoDS5F61P2t0fj/4pd0jWwQEuxyYul
saKY9P4RpmZ5gl9BggWhj0dJs1EQYfrvsDQRtvbx+iZpvCmr6X0qW147lYFoJDwV
H5OVr8b25NukBWDqUpEkrQ/9r/q0YNzxOTzqNIXNxOIFNwU3nSiwE0u0evuurUTD
Sx+lVwPKshLi5mitWQ94YNS7/7SSY5vnukiMf8QFS6GpvsFmpBY120ZNPD5KoyRT
8DSBy2K69+bkE/L4qdr8jnjWkaMK+15BRzGZI+2U7yMOJIComiyVnmISMRk7Eezq
JfwG+1kF/sJJ6DxQjC365VsT8lxXXpJ8jZwgWnRyBo2PYK6QdKIBuchlLzbOPgb7
N2IY7hywQ43kqT1yfg/yr/IC2qF8SbqfnQrko1ctuEhgtO78WpnMCOrJ+GnjVjRO
sJmLjwUWLmuq0to53b6TM3b1Zf8OdfWwgdjIE6Leeepez4HnPeN7tThuYvAybakO
aHQfHjg3BSesUkAYBPfjI4jR1y5TqDdQRZvKtp0jbzgL0R3YEyz/Tg2qnKH1PCyt
yk8Kd+iHblrbGTdhw84XN32F4OGB7piScup9OzkK7yAp1gQ5qW5hUstIz+UYCoIS
PaDVMZsiAxHznHMz5op1sXLcvTKhGybQNqrSol7vuqkhjGUHQ0TYqPyOVDxrAYFl
Z90hD8oMDohGz2e8ZgUYmfFCFUJuonwiB9bdF04cGPNiPZNgSnLdsRhHYnkCIc4O
apDvYUGZtve1rtF6baNdCpjmcFFrbfqZElU/TCF6dqhtvuW08Hg4mOc/xlluViqJ
HjHKMqKRib4/EG24+BdtoBEXqJMYsl2pQTkaSmYNmKtcFwiUglyrmBOH7IVtwh2d
G7uhrr+/XglP81v80po6eFU1SHkG2YK6wdMoR1Auqtz6JL5k/s+PJJD0qgf8RgvE
jIyFemsNZtEus/zs/+ZXdoqPcst1DbQEAUAwmXss+z4mNDzkbGdgI3JDDndLxemB
nUzF7WmeNJWOG+GtC15R3rgxab9dy/o9cZNKf2F+7tChqtjs8uBDkkkXvhgxKvQu
9JwfFRxrvdvmuUFsCyq52sBCwMu91+YW1uQiRd/IscWnSLOCwacqe9EafRhT5kXd
1p8ttFeEZlJToCmTSKJ4eyXiGTfPxD04Y3tX+P5jx/apM7godh6T/s1G3JnvpauE
H8Bc8vDdFbSnJM9XMrl9mn8b9DgPrFyhmmZ6FpaJTjPuAsEPUIGpvJuLKdE1SUk8
LLMm7RhCzCp+NGCauTLDDXY/osBNUdc2GSpVhEKbTwUNuVA/1PDXl16+mfMNH11u
lGgbdSl3EG82HdXOwMpmue91mitN1wnfI2izRY3t7qkMZEhfvaZ4rZhXyHVsoF0O
pbiUbCIjQ89bLUSCuFsljF24h2LN/wWc7WgJTHfKsLw32i+5aoGZZozopjd5GZvJ
zWhE7mY+BFdj1wneKemSgqC7G5O2yAtZX94lV1BjiNqEqlFemiYsvdwcVeZiRIUl
1h7gOvIHk8yXsamq9h0pXO+tN/wVWSSNc19hlR+kIsdBTxLvuDf/sbP342zs04Be
o0LiDKFIa5nnklHl+CmJ/aG0YxHLfG2qdxmuvJS2raKKeJ79IPwiESz3pvYmEAJk
ko0Z4j49qWHBk7ce5AzbN8muKWtqWVRCQBKIkm6JalEuRj5pigVSlKugAE6AoqAT
9gZ8nw8WjehgRPV5EQArHGhuqrRzT/51dZeDkAoVVOlodn4daFxxcqyCB+BiN2uW
fK6BOwB4v1UX9p8DdD3a4cjZP0X2tUD5NKJqypW6DOB/QnqARmLKoqM5tsK6EH5G
nG6f860xDRzXNp2FyrInS3QDARFUvesyFuVm8YF85643kNmqMum2EaoX6frImos8
iilxylAbBhGNeyOz7VGJWexd2Y/gJQznsFcaBkUqxLkeRK4k2NwyN37R6ff9Mheu
2qDRgAYamctOyPTg68aQqfjFoZszbykkqOu18e5X7l4f2rXoGgJDph9JSzB8Nko/
HIBabXiXmcyDYsIJ0uVQLpjUCh0A/MhH1cqclPp+y+zzD4BcFbKgcBSM/G/9jkoB
VP7cnqcKMqwkErSYi6jQbvwqWQ4i24KC6qNDzOd1kYu51Lk/PCjdXFm6NmLQnBBJ
ZzySvi2oPYoOI9KAnrusqMJYwJhMZa82FNwt2i2GTziaUfO47K7feXPydOSjNVgI
0Cp02QcNbPyEvtt5lr2wfRK5CDIFSQ5pPmm2wxqqSQLZ0SxTDECHdZP+suhkRSdx
7Lu5ltfFTZYNldzdRblh1+cMF/Epaqr2KwpSXZ23BGQIGwhgn6tELMBHknuKeTER
HyudENyOiahXfjVMVMJR/61QXTlmg7of8nUk3X1rTBwdr1YGgk1hY/c2QyaD5r+j
iOM1Iw2l2xezX2rOjXDHhzEZVq0H1RDaqfl1T85aaUG9ffdaT77cojmci54g4F6f
GckvUTtFr/hFqOPMPoZec9l+u9PgawGPhfstz2jRb+y9GRLNHvgt5nS5PPokf6w3
VFVu2JA2Z8q35sxNn/lmNLzEF6IsVAWpoDoH9QrB1mEj3m0p/kmTefAlYHxGpsSX
0SfZZC/5ZtGUiIRWI1cDibe0JiBGrHdl+5LoKCXAH1wLWs7kUpK00mAtOEH2nvUF
0GpR29Tf8qRcSLVKgEEqsMRbBZusiEHSt1llGPY3ojopmod0il2zyjEq4spN/uwh
+irP0DN6RKamlUDS6ZlSqCEQpZL7nzQUxKRXYuFs6wNN905q/qLUCD4vfTKyYdJK
V0Znpt8kjRAHL5htGMqIkZTSsnU4cZD5L57OJ65NM1rQ2CSpq/ymgDyxt36s/zo9
OlSHNXuXd6WIRxHzbvXHBfaEJTyt/m4MnvFDfLeW/TpedzIqKhrSSHQEBF66RWJ9
OrlZxhFCg1r2xBS9D28lh5Li3dOh14JRJnkaVwLQUTxoE/NZCfIeA1Ko6uCE5WoK
YTStpV1P7kBuGyWlFWhsBiLV1nsjVZzxykAt5evMhtZ7ca70UMfhfUp+binetazJ
/aeuZEYc4QX7oU0DEbyQCOcbZTajawtlIUWWHIKqFUqEEAiRpoeOz5Cd5D4YnD5b
8SOzt0EOJM4c2Sq3lHg45C0Mk2DCdbGv9HkSENKifkol01K88XuBMYa1OTvFnbdz
HYSetNj31z5pRZx+MUNN7lqooTKkPibObWs6ahg2p+vKSl7FjDApyE9GPRLtmNTE
DpHEAzcIDTqPKnKFrlmzFf3MbX+2y/b9dAAvMiNn+klwVOWWpOBjNEUGHlpTs4kU
LSgVX93gweA3W5sBt/m+Faq51L5lxOE8BM3NUtfK8zK8zzNJN//ii7s+aoloHqhH
z7ol8dksgHqZeTF9OSHZjBea7vrUJb9FMogJ/D3zNfKvwJN5R51JZsSzuh5oXBO3
/ffJKjgZsHv2CfDCt0HMFtRk1I6Z44rtIAfeKyvFkKLoF9QFrua7xQsIRFATIIhV
XYGx4LdQ4Q800J+RSilBGn/mDt+cE+sfv8URxe7lWW1b6nO4eBP+ef7Qi4pP80mc
MHkScBkajiWQiiv0ZfqhoFZG12XHm2Br/T3EiV3g46b1agzR15YXMAydHwlURurI
iubkxI+oZpwojg4U9BQBfz79yDFSOKneOvDA+zWDWYYZWeooz38Su6CuJZVD0TZj
sscgEGmzUnV8sIYkj9mzZrqJsOXu2HwGNSmQgKMqccxS/lpvqwsuL0APbCS6+3S/
A9tJweUFWvcjT+KoiejCqRLeUEFX5GzE6Bb+MZ5pCI17GeKOeNSdvTDhIPYlAzJX
kGKU2h6jnSOI6xmQeds+BvbUHbA0HT0Rqh3CUqyNol2SWm58xOElSPh6bYEKPgaz
P3c3+2aE9V5qfO15w3Y1eCjvozaf7QIjpV5HnhfHuHcMXK7AtStWka40O/gVEc1O
yPVy3Mqulw5s4uNfsNSbPFmiboU21tcNyTCpz9xpGRgHNYmVgr5odklRDpAOPbjj
iTyYfbeCEyRGCAtNrYWTgs0vfaQ0bJ21pv+vrwkCZyCH1/nlbqfHSrgThGVHdW+0
wsPaBcWOTZy+3y0qHyuX6GHcYZXyC3yc738zM/CVMHkQUNHuV+sCqbP9LPADUdPS
KyKOIjgw0T91sdWm0i4Q55990SXOViQ2fCZuBPVk2w9k8wcuVTqecOzxEODoZtXa
BIkePGcUl6inPQ3KeaeyvBu3B2tMSyzXFL0f71w5YXER65WsHDqrIaCthqKXWRK1
2YEli7SQMCQjZoEoxRShk/pnh4Rckai6Sh4fBRG2QgCMzt8FjVH2fQQNm2K/xgUE
F02fOgd9iNSpVBeHndcZdLwH2h1hGD1Ih9okkrECfwORrjyCWvyX2W0wAuvSKtWN
CEyJmDdgpts8ssFIgt7q61VXTK6s/p/5amL6TCdV7YWcPtSu6NRvlOpGiRh4NAND
5NvYcTOq0XkmISxsCc0vDylqs2dqtUI4GAjh7GttWp9gpbWcvI/oJJI8D6pQSKex
HWE++PU8biLSKJfirHqkkPjw6lSRLiEpE6iNBxPajLkbCJFMnrnuKpWsTaXP80Qn
o/a3Dw/bC4J5X/fIbY61TNdXLnNrrH+mAYRq2hTK39p45BxEuN8pbTr64jVRG4Sf
AByrhC0fwPcXxgJ60U72mh0TXYydIORQpIDACI6TdKlM7Zk4yfbo+wVYrvT1Rfv7
u4n2/A1MjZTRIiRbjD7DGQp3ATS1akZQ7KByrbGegl0HrTudvY1lw8ZDPSgnPcTv
qMRxZxjGAVg8SFAKkbjHD1+71Xtg5pqR4mwt/6HlgG82sbdKa98lz7QpFcV63QB0
fZJ5fs95lOCzLrcDT70JrleyaCq9a4Y275rXpkAlAI5RVy3uu9BOe4AAH4DymLld
G4x4tOqrzTUN5fhZims1KT/U4KBvMRT58442XiCNZQLGHPS+h3941t52ouL9YMKM
MMu8YhykZFQrawNydmbbZ/vF3w8GuuhuKwbBvpvJtjmxzHjZClkqekKX7LLmZSYE
tHCv8Un10Z9i/IGoHj9RoX1lZXxsj/WOiq5CdhFkcyHbIy50OkaLMEWNOkyWQYRu
fWvhkdIBWV3qRIgr7xijbIw6BQqedHOMa0SRqk8tAMwaOWuf5K8dBKRNwS31RYD6
7saJxAw5RZR3apuunjRPMx6OoaMIdLgCGp5v/GbQ7lkyKPQlM3kldOXtJ0BJCNlO
rSwNAQTuay4ksl4iLJBqgKA8l4XU1ZLE0faxjhaTD6WoWjk2Gx8zqEP9FIFhvkMz
cIKY8M04edCLzP8PNMkN5byu0Mw7M1CCtseAgutYC65BRlkZFvWL8Id0hDW5JdPU
SLhkVg/tq0+ImchTwfuwhsAdJ7eZbV8MkCUB736tQlZ7nrQPCNnpfqQKwK5gZbml
g4D6GcxNvh/gWb0EFiNh5p9iOexjIRiioR7Nsg2J7fTyo7vGmfK+QcG6UIYcFlpx
lFHSdPbbhucm2jRrPK3ILP3lDjrZXlqGEiMsPI0b8nCJ997CJN5rrTpkPeHToH6+
aIfhr+Nm3tlAOBhEnRYEtv3nmHjvzu5lXffOCqyn+t7HAXQwdBuwHqXUWU0P44es
cNV7QnqMjKyLxHJ19ssuUg69Zt2H1pvYgA/8mJvqslXMVx9s69tlRbjtfpk9aUgh
ZMvx28+evQ2ezWCJcQr1OJZIZOLvMhBvEucA1jIb6F+Rg6ssGlVkFj1lBJ3RB9W1
qYJVcATwY5QEfoVp0A39XPxg4ZW+3Jg6qBAO3uB1skCpagp0XINKThxWk8Wn8LpB
ySFYYXTRigvjp/OQFVxpUTEThbeq9GdGUrqQr/YcNoPwjarmy8WCTHdywSejlcmU
FUWWfMxH5aG2Q3nw0MTcXBR5Fqn2nCAB2kzo5cPYXs57Nj9kNIcbAWJNL7bSzo0Z
LTSJ8Y+rTeQpo0xLQTjjeH/M2LDVfaCKsJKwTDJCaMqOTZZ/wQqbJQApD7pxVrNL
fwfEzMbXNnKeTp26MWz0d1TqsAj28P1FEewabLKogqusz0zW6aaSxXJjujaEAROp
FaVpcg/tIGCJm0EJwONGoodecsPtA3VhAg4Q1M7DkKNC1zDtUPFi/dqZkw/td8Ih
OaO4AutUSg7obW6FsvRCQvwQinzXcwsYtAS5BTQ735a109TeWRh4jbboR37CrH1H
94TNgwrvBKOzvHrK/Pr3D1DIcuxswkOLmPfCZawMs87xlmyIHMUYFCCK8tetIpGT
lsncFmUC1TDFXDQmxCcp4yLSPKKePHldA4GePABkDzVaYaCHddjac2/pDho0G6Db
0XXb2RCKIwayCBxo158qpLzrabX4yYuUOnukPzVl2od3jfCk4ld9YvZ/FUA3PrCL
agiumg0hbMXN1qJ2Bc6HmKJsW0WqDaYYk+MeO1eAExbJTiYnFfypc5P4zBA0eHPj
vkhIFst1JKhwmeUbOumT4pAY5+LGufO/TUrGv1hkfxSHTY3dz7IVFyETsvwdM6OJ
VzHJ/0JyXC/NFjtZopZ7ORoRo6O3WxqOFxoydvklbMQtsqW4i2EpHz2TtwO8s8Nz
Uq9FhtR9qERFRJrNGVBjBUj/qCgZMv70tIcDmb37aVzmH5L1rEReOR7WxBzg1VRk
kNQB+980bJznhWCqmjj+hTG6xx4Td5SCo74aY3AXNNhIkMeRNqEvNowPh8ikOnqO
F80iT40BLpvfrHhp8ZNCSEGhM89bvUEejyfewlNfUhutlrQmbS/YfPnZaozaJnSi
93dqp4YDdGZUn3n5D/YXEbgytjwcorEPKqRkVJaRref5RYx7XcW6JSD5BC5jBi5o
I96SuXBQLn8SHtri3g2QPk6grDozxBbjoAyGApLS4Qa9DCcgW2MSOtv8vxrpE8IH
PB2ljruQfuqTgkLiXZpycK0j+cpLHrnQROxmEqFvuqaIXrodMHYvOVIPwQIHTEvh
0+dcQg3iL52L72Rxa9uWS0fcH9ZJ37LYv1gyKdHKiWLiC9WuG3q9dRgqVfoPaSoF
Ihizsz+O/Y6QWrl9cfO5PcpJvBvgyhtR001o+B9MSal9iSoYqeqccjFtoLtzZLEV
77CY+nEvy053cJ+QdF+Bb5aztBnklAKgZ4fp1XgubGPYFYNUwcXNOUxxLe2Tv+Fg
AkG63QLxyN1yrzs05PP37kPo5BWaN70gzOZvhPBjvdy+B8JzwKHA/wCYW6UMrXk8
yWtHzeZ+KlAGengwwpIWMo14/3/uLEF70siWVqne0dA9HRshdkNP5g4RZPtAdBld
1n/hVbN1A7QKa/C6lXg0VcHGZpwVmE/4v3yu1ZoDz+yZfTBQ+Pe87OO0XU87Hk1r
9qHrDaLRDYNOdZTOz0iL0/9VVEYwyzPI7odD++Dbi9D2hof93ZXrWGd72mQdJP00
o55dH6o6bYuU6E64ds7BGPFXbPed8VrjCZ/mz4PiLb7l4s0vF0mNiXIImUvQ/avx
/tIS4fsGq6FXWBL/ZsJpHKqF+OqOPvvUawXfkk8UOVW+NRMambTAH0/dFwNekLfZ
/viUVrOOZTB/WQeAAlTnnANyQzjN8cRNCsXHkLMMWFM89nflCVLfXwON5SOIPP8+
vxpUA6JdPcpUrenPWnfXPSlqczLBhLlhrarxGnQa8MaD/id0+/y7qqbQMXtNXk8N
h3s0zCu2Gn8gt3YumaLyNKBGR23c2bXesPr6v1f2TCoL77r5Dw8djWp6stFMQ5zW
y+TbvvHtbPsWqz3sIQWh43g/6klqTi41qft8qUPDvIcvhP8chVP5Y+nhpNZUFWCj
XbybPZw9YtAJCa/kfkRjdl1BAOmWWG3fWuB/eiEKEVXXuk3vF64i62Ll0OcktlFC
LAsED3ZQcWSElZrTxgOuR48c0Bv4ATvGVfdUE0/7Ak4IqQvDTLJpSVS/JUeZus6l
vXw5g3kKKQWbzj6+9xToC+93BRV+jNePxZQgQ2up5dc1NNtTgWOA+hJSNrEhZfb3
eh3VMYxDIRtPguhP2NyCu0Zip0vRvneu6WaCcSyMzG+lqz16Ry8TWLoNmX7nxukk
G6EvWwoIJyItQFq7wYxgEOSOBc67mVbHAP1mwwVECmmfPJCXvjkEvmTZjdtfZecR
2fzZBNyFVKUin+2EVsbL5rcboHnc6oMidq2+7aMFv7Ln32iweW2Y20eJM9OfX7Qx
pdu5qKC2SJZE1csTiLzT/iHKA+ccjhQWU86cIAIlWhuHgnOyDi/wzRD6TSrKXMvP
7NYAAuKFn4DK0NLt1T1i+cYIFpBIIC8cjCN2LJ8r1VnyOHly8Z4vfezukpaWVLMQ
Ni323Ig40Cnc3di7Wn96TfU/PyK25JSi4ECKdU3DsszTIDDkdv1pZrttzOCAm143
+OSNVmfygCOA4oBIpFvEmmhvVEQ0I3KqYxuEt8EXSb1QIWfIqpM5TvodEPaARch/
Anz9sLWnBlNo1fb+9aWwyreHeztmDzrWSsUu7cgvhJ5PIeYsoKbYsHLRebn1E9jS
nvZqDtWX5OtkrqV6TbqP/VxE+D6AVmCC1BCZlQN6EYByspVp+kDrTFBJycbHhnq3
VrJUbDaJkqAcCoC3jjwpuNnmG3dwMMC2jJ8tMRV1CeVwHAWt5LfrHvItZ9uh4qKN
zsTXwN3HDnBjlPfCiGFC9yZL61xLKH1DU4+7JySDINiVQulRKu75J5hNr6btk3ZR
CoZyJ0zv+JmK0Zg4p215kuLl1BPH1k4iNRhpjdfiDUKjI6mDPwpuP8oG55afFb/a
r9tsKLY+nvKTk2wUzj5/TD++BoX0j/WhBhEWSeVCH+PUTGTErxJLWkApeLHxSeSf
/607aBip2gGQ7oNVxuEJC7gXsMnz99SGkot9tF8EOXPPYZj/W8CLUDhysu0DLDTa
CnQGiWlzxPm77Tsy9DQHONIVIm4ljPWKVhfaBL+ws4KJ1tKGEfoUEBH2bNs91ZCo
2ie3f+uYWcVFZLFMZGSI9hGNu5mqPKxnyR1LMaTPZJnfRdrDnAQxXteHz+nni9lk
3ZXgVjFYslkZ346VvX1H02BSR6mH6y+Xpx/bdp0Pb1RfmksP5KSzGGL4ASCsK59G
JzPVFDHvlpnkVeTCHKFuWESBJBhHK9i5IWRdAxwVAXFnpfXNk3Rh7QZ33qaqlwYk
bXkjTv0pFeaUYrD6DzpvsyP6vS2oy6GHibESeYpEdpb2x35llN+tScoPCEDO/xt0
nifRr2u3NN2WnaxzxmvCUJl3WX+6+/3+kfAOcxVlwyOTRR9ymvy02aIOV0nITMY+
EBuel2JWKH7Xzv8evyD5ibvHaMVBL90skSiHz328XujdsDCoF1HPyRMgYfOekPLG
08+H641OB8fYD02f6ei4bhMkVBKGlKHHT/82SfnK+oh+KfVr8Cg4/CSCf2i/Je0Y
Gle+Da18H1sG8l9C8JOsIOt5pBx86EqQIoVWWGwU/E2HBt97NkMdud5JIxYJWAgJ
pLdPFOuzl7wNzGzHhzvc6uSNBgyQa+TgtgueUQWslt5yFmgHEm8MdNPiySHsK1BE
1Rq2fssyyJGYo+xX4ipQUc7fi3CrFx7cndRjJpT7BaZLUo/sG6YVtjM3QgSDnjun
nxeFCASeJzQEisFlUjRPBtVEVsaJUArVg/dR4Rkf3n2HP16N2b43mu9mJ+50Ev1f
YZ7bFLnTW6iXZzDcHToDRxcxj5iQ8qJdHlWTOZEpnSF+ShWgwORH6vcmTT4ygwND
JSghJ+53m9QIymZc58unRM13/CNRuPW0iDKuYRuECGlok7wfhip/2EPfQMNJj5eF
`pragma protect end_protected
