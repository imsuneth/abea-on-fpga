// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bOSSf60Gw0CmfGFYjIccQIz1PbRPB2vh72K7RMZc/PjJmLZS2MG1LkSPQbIYADoG
tD5aakhjlMZkvovLz2vNdMhk3ziOXSWNV6gabG5/0uT4lnfLJQRM9cosOynNV1jU
EuZF3wUfQt/wo1wkGvmdaOwucNd7V0Xf1bh6ttQxAEo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4016)
SMOgzOvepfdGtfi+ES+4K7NaXEAgkf5c4El/qqJVw+WC3EqtkadT5TtMULcz4R17
MksL8PG0r/N1mtpWrJjxOwoS/qSaMIA7bmU6cFGr0jxOjS+G/Tg4k63TY/qKRJw2
CSLjRAkWDxMfzRWHVE8hzOM/3On1WfI77rTx2qlxD6KCnbRBjc3BhnA1WZUCtqo1
ZTt4FMJJ2xlz5xsEgSRYhz9pMw/CJHav6lf09egPL3JgWcJWwOmmaB4No33q0vfY
XjNtYWrpvCxmoJRyv1I2K27YKeN1Iyuf4E9tbLMEq97cMRLDPjWyC4S7m52eTzGn
yX+r0vIbqlPxI5bqCO340bITSCbbqP6vb6BgqwRjQ7v3PMtPCFMSrl5hv6YRqLMc
voAevpC5BAwgrF57dF1Gqu3Mn8/eYBMbbksbSKffOhZZHJkjXCxlQUouKDvJw4LR
R6k4TvshyW2UQJdj5/0WyxuYP3PBqckXiLaKWCn2hznPey4qEHseKmNixCJoBUa4
htNxFav0umw2biZaa00x/E5kpukYZsZRcHQvRNvR04Q7Pue/vHokEpfeM45onswZ
wcbReuZQu5rkoX1Jp6qtbDS4MXjN1CtVWGIuT3ys0x6kujqNxtPkbh87MSYNHiRc
TomN9k7XyKinJBBkE2A6D+7uqM+mDV9rSE5r4dQQFK6RjIp1sp/MDVh8ckFjA08R
BIC7TToEtR/SWuKSnOsQCzfYojlBHHO+Uft73gmv/6y8W94nuUUcXgQXu+wrl8R4
0tt5tiBHOT1aGvo1700p1ljhHzCBa9U9mesXX1SHAz6wcx9/3SzRm0wNSW6cTTbP
4Mc9xNPQ5d2nrE8e5thqZqiTA6maMPUL+DTMNhG8BBv1M6wgUoUtxiReOR9AGva4
H3xExYCUWlCxSpXatTjV+A5xnGhyDxD3raEJvRsOAU0d/hPwtRAfa6PUej+lzRqa
Hxy1o+kWqa4EkpQHy6DjCY4kaYCk7X6DSgbqY6Fo/0gOx/ASfB8uL2yO0bWQVtXp
eM6kJi7QDlEPSYAPPtY+JZ7Vms8oI2UUkktx8WmHhC8CIaGplbSzk5kSMID7SdAL
78US9mb4n8FWl65DGquiDSrKlepcdXdSr6l+9chQ9XZqZ+YW4oSGZk+7UjRS50le
PstduU9wPf4CrQovNE8YUER++q5uhKreSxsrtQO/A2BYaSVTynZPkFkzxeWTNbMu
99rH0mOdrgY3uvJa0JF+wI6G1dH+oT4y1m+fgIANIiyQHZ0T6JgruYnLRH0IFRc4
cCvAQqv713V8Jkeekw9bk1jSM/2lXhwSFrk9ytoHzF53hKzR3VaJAY+WWYORgWvl
u32sJWuyPL25+3vu/9U7zrlaZECJrvX4FGJpAwzYFFJIgHr/GFq4qgGIA1VnF+Wr
9qeMN9mXQoioDIzKNOrIrwm2TORlGQDVk4M6m/SpF9PKuhx03yh+r5D3dHlHz1Bq
5dExXZvHtOSSpGd/V6/BIs3ETtd73kmR2qk65bR3dpFKbvf2w2StIeOQeqLjDD3w
wHn+wE5jDHgK2CsrmmVsf40V8/JIdM1TpSoBu8J3bsANDHsf9XbchVND9ESKnuUM
7d3vqZCRFdlDZzSzzs2J2uP23pZ5kVI1iwI2ihRRgPZA1ZHdXcjjlMGC5DoDD9RX
UEUt41lA1yjGRLa+YsqZuAmvf+xzGooDGwFSHfkA61CKm1VV5NwXF9pxr0Qnzd5j
lkOM1Jqk6gFVM/H3VKpfcQCX4IHFiUBtAVY7azJ6PR/JTUD9XcYYaPWR4zCmTHiZ
NB0J5jzjZQf0HufvtU+kpcPP2Fb4u4WZDVPdSJ91qfUEDFJ8UyDgBYIJ9Dk0bNoc
o+ETFg8EztZTYcnLnqalSwfq7bsaUCO1ZiNg82PMGdDf55lJFDohJX1WQVKPPht8
HvSZ8OOdK358jYlwFIYUieNmH0FHjhUqIZGln6wVXfBtm8W40t55hDXIjAHf/FPW
RcAD1jRvqXkKC+lvZKH1UJL8t2mrQovR7rUJu9ohEtH2k7GQu8l198Zoj07MYxpC
nzc/y+Ch688puTTXQABcbWE3+JuU9oaBq6sdGLoEsgOcbGUi4n3Xk5iZxKg5zSqZ
QuDX2JXxKQBq6FTD1rG0QKNoSa2hMpe6CwNaTPu7uFT791Mttk0wKaJnLlPUvP7/
Y/YZSboJWBEkBE2cE7W49mdfmwv5NCsbWOh6Yr0GvjQTERGjRntfFbZo84GaDwwP
ftZZjBjQgbhdtxPpcSOEqC/SPaCGJ+szijhz/UMb2eaje/jSKhBHUDukwS5IcT/B
PRIoCNf3v5EndmPac/bXHYYI1XIvosqBeq02kicmOBupscTPVRPQlJ9rzlReAs0v
iSHvYYPZuP1xgD3CVsciogZuguwHlYQWkdqWUwzgaWkwBYleAM6G+fv+oPA9c7D2
OvEq68m7ZnzBizMb1RS+4jbYD6e3LNUSRNeQYfPcA+0XQhfYAc6DbmxE0ehfjdfI
d8x88RNCFpcQoKf5o11+YyYUqkMOReeGano97UTM9wXaKT79d/ccWYUxQRp1KRJE
QEsH683FDil8eMQ/M0BqxbPRaCPtgbgYqrTdf5iRnrLdltRRpKSnjwArEeruhgcl
zrX0PWm6nfAY/Tu5fUzI8p3DEbzNM2cqpCmMPbJIb0cHOZjKkpWSAsayCK6FDl5D
X2cEim5D8tv2OTl9/eLcO/TYzqL7sBHw5xFJc/SUSJnoqiC6K4gTD2uQtEgwNLZO
9RjqmbLqguRlVMM2ZLo4rmxvqaKwjwOBHGF3EraxZUK99J8+pIVmpE8jbnSiWSnh
pWZiTVFmo1A2kL39WDif9NmkcWYqfCsBeHJPVfQFTFX972JjFQ4P5MsoKN7UsOKX
BnSOGFZIt0J4qm2S8IeEZ+C8WUjZPVg+MZ+7ZKd/9ECIjXgnvOUMPWkc0nFTHBUo
UmOWKVV2BH8T21GVyXu+Wn94buSXx4UTMcL710eVCwSZUi6ZS7R4dwJSugoJq5yD
3Sd8p2xzSlDDWy8tRGj2RfYMkurqQc0eSDinJYxXcosy074EEi+n+LLDvM0e83cI
6AlzWd6Ry5fuDC8UgfliJWypBLd+JFfpYLNBbFxU29tqoUNgwg3+FSThPJOaz7rx
0Q4GWEvtOqvuR90Fukfcn6B7SM5ym/uT8U3KoIjIOaH2mqtPrF1JuRXdk+PDZdyf
PShuqEGHpyQf7N1fcPaYBZWGbj5yjV4wX53pt4aS9a13JXpZ6C1Q9qDPEP73AIkx
1Bfp01Zp/DE1zZF4NM+EH6wCea7SgNHOc5gaz0TL5s6xqB7QJ9av+z0dcCcZbMAx
c6C3w63FLH0ql6EEEzu2dvMOIf5L3PvjVGWHyoEmxvm7R7oDjwjZKXPUUxPwVDc0
yg3kf4OSEhS4tCn2pWGeo9q+g1vi8/5HveI9RZ+7tPbFYfZcgE9RNyUdbclNsZwf
wV1iA0RgESrIiXNJal9Lar+XLwKTg/FylmZq09H/E3hhzU/50pSvUwFdK82jmIlj
6MC46SeIg1L8MUrxZDBk1ekoI4yv+wWoVC3WZCxX8ZfjbUS06QScltFDPXA8oVhN
yUPttg5DnlfLAXpnw9rPItWwSBkgGg8FJjOCoaFzNxl6SNOnLNKIlkIzLjI69Smh
xtqNv7fxKUtYcjYG5eYH4m2qeuafs3N5BWFrteDhMiS0DvDaET1wbQxHXT9nBE3O
o3UvXgLO2KVajlox8wOJQKSatukjYUhX47AnYlEBXPJQETyX975oKgo5ZhjF9/8h
Kn1Ztx8en6PyMeVSQgzcvkxu9VW64LaJ1U9j3B3QpdK6cd460AihG7AIJiCZaq56
UxWfbEIEJSr9H+Bw3EIpSBI7H+Fbedu4n/lBu4Ovh3gK5K5o7jiIRTiHHYjQuM/+
Bl/0LJhFoiQ7DCSRzS0pshXW7zzFEP8tmBbZhkMdUb17U6JxMOEW1oYMLxlL12IV
bqX0LzLuqD/p7VIEUOEXOKC+yKz0xEKM4RAiU1Ca6pk2ONTnligjyOwU13VswvMO
tMCoU3Czk98OjLeYi88gqQGOCQu04rBVO4ZiZ2jMKHaaQGy3KmJ4oKYk32DP9k+l
r+La6N997CEfhaoFvtXi06NJKyOfyBl4hYmChZntgatFG+cHiUY6oYXaEzeUVgT9
7tWS2RgwE4nOUjMKmCSPXCVGgsSWGNpITTQsh/4fWjUpGTGTKc+pVP9B+wxMQBFT
MuBX9T2iax+ueL9ScL58ZMaD2d7NbPPBOwwkTrYzK5+pB4fwPZQZIpYHlwwHEC4x
C1e4FWUsjGMWumZvnaA8+XemqwcqFj5AxrkrMt69PFWkBdmZTJSQZDdcxK/4PYpQ
3drnXhEKSJlnmdcQ3k6jol/zGBXR/xDDZ/LknOQWWwBNnX6BD5AiH3Jr+lfE1xhq
pShF95SQwWk5ovp0Jsrm0KZ2CWPAEl6eenLjcTaQpF8NVgDT2OnEaPk0E9isXLAp
aS4SGDrTRjkCnN+K8B2D2YGQT6L+zzXDfsHtf0H/aUR3sb5MmzargGgEVZ9ukdjp
fxmLgNqOq1/y9N6HhsQjPN/fSxInWOWjWulL/2MJcNwzicegFWZOQUWq5SyNs3hz
FmjshEeewCBtPjgIpoyAbKwr37UHbNFzUZOeJaR7uQgvSQV9YOIiEiMXqsb58iKx
2AJ0QZWKTiJrBHsqyoP11FTrpM+C5xBAQgyUsmx48OeAbd9hYA3fudjuUZPoSqDk
ZmqHGrTvwpkIMC75v2jDClwxkAxJw+bgsykXy7g52ZMm4v3kqWz44xTuDUaKCwEr
fC92TN2lBTt36o9QLtp22W0jhyY32rJlYTxHV+xUZMBhPHrN0Jw/8lCKNDd+CrrI
nE4d/OUgmdZe7jWenphiIOgLakBwSeJhulSLUz90q2CkHuwx7KONyLSnQfHSaJra
4e9uY6CVgM11uKtv4O6MtuyQSF7BwiCwRWyIUqG1OHr7xCnykxg9kZxZP2C0rr2P
kWnUGmsQ7kPuSbk8S/CTA1B7fTYsBPa7j97F4Nt+X8vrEBe41EhoOnruhD/02pdU
IPFRcczLKtzN7MsnqyxeeR7qZ8OqBPIYx5WugpORfxxfUTfCWg61MbjY57Z4skEA
HNYXOMNV22oDgLT39Iws6KfR6Py8SEt3pkOVjkj/Uo2ceGVIXIMuMwYl0h+7P46F
XQ2H9mF7mD43d4iwFso0f5BzuIEnBLVTtEbBrLub12UlHbBUAwdyP8ORtr5jDVe/
ekN/2L4djT15F/ucKuejPqoOv2dPU/jd0a8GBLl+b5DfalYrqbwd4nHAKLC4ReFx
DXKmcMe/oORh/R8gyJfqUTe2xb4paoa86vyjWB1DA+Y=
`pragma protect end_protected
