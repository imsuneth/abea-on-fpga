// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:29 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LcYwidSadz3oskJ2Ij0JBouDvNkB+NOOfxVb6v1Yu2o1OCZsn2H74BNMR8EXZoR0
xPEJk/3jDuUvxSV2v+wcY9eZa59MBGztO8IBL3Yr/6hXGyJCQvVuIySokvQcPRoK
xN4zOKa8/QbWe3Xa8SnzgIQGrv4Pb9uaTn1QPsty568=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46192)
5DHLzSnWHdka24u8KQuU06hFob5VmFwFUO4s6T3s4Ms+bQ1Sm5JDJ6Zq5qCM5GP5
2ni1sqAjhXX3n2EpB7gg9o2tpPG4Zm9Jep8cjt4XJyFK3/HmiyMoUboL+NNOmedv
D0pvNx/aRxzlMJ+hqrPQ1xpE2V7he2RDQN9Dn4lfL4zouyPlbe0B2/u2kWvmrDDx
pTr0vMevsiPey8cP0ix7BP9rpJXGR9wf3xz0AR/vHOQuSF9g4mejDI7Cn29jd3vP
RVz72RgMVewpc0+Z55jU6KFf4jhMp1uN7UYtkMGGhtEI4cg4Dem/4tOTwannJYth
LlXG6FXZTwuoNL0qFNEq2b6bkY+VT6IeGoQYBg4eRXEvTudEFFkZt9RFhki4Czuq
qikXlzV/Mh5yzM6bMilH/TZm/h4a40hnqGwnZGvuH7HJ5oavniooLl7K+6IMDZnx
Yc2Dg0Ez90apbMyH8qkt0Q8LqF1co/VuMhY9vrO2RMEYo+kdWu3SB1rRWZRzZNq/
zcyQhINcqg/NutDdSxHJFUI4u9YO0a9wwCnt8NbXC/FWPqomojRztNSyNH0PqcrN
sattKJCDX3W6vMbBfO8zd/2BZH+AdXXQqBvGQjXWGqmjkgnrY3zsks1mBPN1rfQ6
jT2WQOzqto5pO2E9SYPZ45Oo7zgH12dy4JIpTY9z0E3i+4kkkJ9JHrvYjKgEiAHF
J77gFRsUsezzgtrJCkWipFAJmBzwlnEknGyWnu84lrdAD+Cfb8e1cbrjECSG8OeF
jqGIJ6fmt0pQOLxUp++z4cQrnJqmLnwHlFpcLff16nSWE8wm1FpKnmPdizLkd+1F
xMJOcnbLRlOedZ2mwRPDygju+WhNa92u52oIj40g2H18NDgUnNBb7qQ6vI/cqOCF
f0tZUAE9J1uD520w7JiyTeYIdIuLak1F9j9AvqfXoUtOGE9uDT5zFPGyXsTpVbEY
uDlpd9+HyklIlY7IDBzywSn7OBoN+el95ijVFy11XVWCzIPWFKLJ7kPk02BUxnBP
QLqALFwAVzm42K9K60NNK0e7/2z1jeqGaz6y70CY7Ab66OWUB0aJ0up7u+iP8/VR
OdgjAtIw2ziS/VyyIFuDiPeo8pijPDBRV+iYrBvt52955oRfqPUB6etdqj0zrHEn
gLaDSAYUWKXbchR/D7mHFZ4CB8KeWY7887eIXHAijSzE1sQl0+TQBUnFIfgpFAcw
qo/+jiG0knYVXd0BHW/YakkvVY4hEUgyD7BizOntwjazoVDSD0WafMc7roWfYiPE
S396iwCS0Du4Sak6dTITAzyrj/fKPzNneKyoaP5r5llsDF1N+6GDlFuCbmN1AAIv
XM7H2deZNtNXJbRbqptCLUPgmUINLX9xGJ2bE5bepzyYbHB5Ggx7MOvX1Nj1JTTs
j8+YZkNoTQR8EoelXuKXEWUJcezNmfb6VeYswJ9FkBkKGyvraUH7jBNl9ZDmFfe1
IZD+lyVnFb9UILVxbPRDgJDOOxXQBkPBhUgpiL+9yoof7jfyTBdAW5KbBZyOGDkt
cPJFTKI/4kIscpQkIVsoBK1DmG7z2Fh7fEnfTCyuH16iR+KytjMeQc4p0amKUuzh
q04WgLzrfKhMJGku0VmAGmw0SaDrMIstv3LcMj2pTjiwojaQ6PILQYQqnzecx72X
nsClqac+bsnJ5XQCuZ+WxLhLPy2C2vDvbLricRNcdamM6yv0BVtdRVhaGIApdw7h
JHViV8Y+mTCo4us/zjJHbxQb6CBccPLfJBOCp2MqcWDIhzRj7TJQgM///NYuZIAf
mLotstV0y8L/DGhmT2ehnjQ9ojl5kSeTzBCrR0UckY8Px7AmUs587r7CRwzW1flk
qVLFkmp/03NqlLGtRVGggsT6uu/5Xv5dd84DlsRCz3q7PMrtm3cvt+ZkHg3/0jDz
8ooCG7oSvN3r/5Q3VcaF1Qphb2zOZsDhENr/YvQ+Vh0eu0WNb+QlxhPs2b1N2bLs
1+xuQ6zZNPJOkd7C284yB/ZhMCd9TsGj+GjFKvFgtmAze8nDFN+c8egsKMVtPdvd
l1todaZWRBHavqp5ApFV9jPBQQd+jVMxvozb7K78jH2gG/kukO9JuT/xqb2D63sy
RaInUK9sboI2Sx4BGzfh0GSWPprHf9d6uHGBru24JKpBz83iDop/xMaEuSXrzF72
pDG4tbiLY/2NFX2hlenwlo1xpA+Uqd9r3yC21uorqtxKbUmVUHPe8z7ILyNdbG2s
NpT9pzKIqqzmazh7mSntx6EZEvFHsWx+f6d9JWPiuR15Dkk2XeYBmkh5nuT/8cIQ
+6dUOj0CX1QY7DSry81LNVxss8gN1hZPNV2JxDrh2bxsydmpOvs2fSTH1AvAGlEz
vuP3w7wjSzToVRXHaeREmAkG/skLfOkoTPoHrayCbdAiYrGuT6f3nUrETcRHQF+w
sQHVwewpNQnR/DKAcPdDpIdDcl068XvhTU+7MOp0ZclWE8wPI1+4eM+/wOcKefNt
SYdPXkAik0NSlt30dIwbPjJA9PsMLykoN3x7lJ/jBOxyGxs9PGEeWhAS+n61++SW
6j1932CoGNmwywmo08doq8EoUCWrpo1EkcZkZa2WuVe9+zP2rW1BQNOuPwVHTdq3
aAkN5X7tVm952vy1FGXm/Z0vPQUPw1nY2I2+a9cxS6kMHPnCD62TRItuKtwhV2+L
iioGB6oIvZ+gLRSj2qjxGW/8C9JWVRZqX/ohFsSsPS+26GNToo+X7BCoItDx3npC
Sj0YAZnpLbeHvaYqK3tPTr1npRxpJ72iftg8vAAiSiav/BWL4Ujqq82/ygOZ04Cw
wXutLQGXa9KMOz2LUpRRgUUR2kak8Ucrl62Ek7E8/fTLolN70Gqxqrw8vUYR5O9r
fIhvOc6wNFRs/DmvwT3Hvf8erNWrvX7MnUp+jePr+dYrBBaYyWnOXkYVL4LzOkx7
VWP8iksbMkctcIrcMm7vIdvQE4o1hcjvs0X7OqQoQRm8J8iQETNoMhSJ7cPIq/4l
/nzcYo77sQ9QGAsDX05ZZKs8G9hroxVx8knAJSETeEm1RtKsUxCiB1jjNnJUq5OJ
JCJ5OMIo4Ft26Y+f2FjB/iI+JjTMxLeVUS6UVpz5DrfGzkn+9djytlIyNESeoTuo
8Xwu0wn9hO0jYGuY6IXV6GfsByTfmTbY9E9C56yx32IjKIi3WTLGxADDkS6WvEWF
8x0rwZtDFMMWe8TLEj32VxfwoXTfNAO6uYAz8JgnLfuCjRdUoMS+FHPsyBRpQzH0
WEPOwIhK5Zo3/RsncSlWwkFie409pPJXiIBx1Ji/daURi8J86iVKDwGVONy4rlEl
n9wFQ8ia03xKOhfPrIUKcalKcKsLgi7GgzO09vBjLL4GGfNK6T7Pyd1WUoKzVN2q
2K4UXD3JMk5vVqrK4z/5qX+i9YtOqwujZuZeVKXjJ82FBxdaFLDihISYUKRoUicH
1d8lyONji5HElQZGNKZketci55JfzeUfyX0Xw6wHhza4C0ReL4x7mt8LUIJsg8UU
7LnynwKJdOa9SiV/VeIEEax3hWkZo7HTyHFHWAStwkLjDkuNlpSjq6oX7XV7P/XM
7513Ij491nzH9rgBJbl7P6PwoIiULUczrtlLvu+ta9bNEuT8+AkWVAiya8Vp7Sfr
bcLf+m0lAaWzCeuQz0cnjZtxZHNSjyumcLDukG9m3MbY9o3lvjyqvzrCadj3m30b
NQKE/dW8XwJOBqxU9Rd4p9hM3ywt+k4jR1Czz5oMJkdJZyc6+9sY9Dasp9JdQMxT
uOZiUI/JMNh4kh/9EhJyLPIrnSSW54p3y8quidTwhTiNmZIeuBa/oQaguP7sCW1Z
UfnrCYAPXxXcU3el1pKdBku8Yl8JMjqYJhFRAO18ZlXKJ2ecJ7N/elno0O9PjG0g
lbX7e//N6PpprAQOrCqXHzWxDLwtOzi/idtg5R/wpeqyBY8imkXMP1NfcuP8gxEB
VEgUmH+3gpyilNEGfPEpnn+DGwuBq24w0ZTwcD6sadQct72qQURnP0JnnPW3GTld
Z0cFzRent94euEg1dVwQW2WqUDSLTPzm+l/3a292jfUpRh3ZRAuuYNU4I4U7oXHh
1n0OkUte0CAeaU/rlYGalQR9VZN3K33oaI398UiIa53W1AJb726G47jv3ows1ZfF
FruLsgjv9ne8chukrqWb+Uf1uamo7FfCcOiiIqAQ5Ok/XQQouCmoc6Y98qIORg6H
OQ6ihH2zCZEvIYRd8P8AuMr8x/CienjnJsO3P9Q9dBozxBG3qzirQCIJtLzoxEVc
s0OTYYx5CviAtU9x/4gPvD2uKwzK0XBDId5gmrIsg6AAoWhGztFTlhU8XRGwuAfL
O0KQR5+xOPASIRhzbfVJE6Nwez8VYkdem7F6Rg9MVUnV/UKezqIYPuuO6Z6j6dPg
mvEox9IvROhxqc2TTEhCjhzEwK+8aj2TrdYVbzcT4xThi8ZIFA8maY85tmzPM1Bs
GNc8j9Y3/GAcdSGenXhOOKhcZtsS4FgSBJPNdWuu9g6vtX/ks5asMPOefYF+rag0
9Xpz+DY8h1A0aXwKRS9sp6IWB3cHJTofFE4LFSUXhIj4coVoBNnBbLeDDrhM1Jqe
V7Re2jdTHJdThn2J5gLiGZeVrOkDLDAq0Zjsy+M8mpXMNzE8dWP0P04Pm6uIxUhF
7D/6Tislgji+1XHypkyCNU3UIImOxpCWAC6gLhwUIZUtVhqfcJfr/s0UX53toCmG
J3NqBVHAnBJZ1zjM6p6SpBC94xwNUX1OCPVbkZZnxOzAJvYyDiOoLEl46Q36tBBX
Rp6ZW8zC1HAzFnrUaBvQrYOToDp0UV+X/Pbeg1d486qCGwAwIiBZC/fcX5+WxZye
i+bazO12MOk23apxS+jPWO/1QSbYMDmqlgAZbR82atv9L9zA6a2qWKha0m04L+BX
p+9vtAcoCE8m+YHw0eHG5nJGTtTqnjm/PYxgkAXoG4ODZ+f1z2Xu+dxD+fJp0xn5
4k7BPCvxVdDeKQVOMFg6tB8r22/TBUFX+E0UTK8DD8IK5AFxKaPaanX8vHCXy6FF
rALesedvDIcPWlod/2MCZRB4w1SFPXpyT+JiVeAkiHkZh/+lnPSpX5xwuqq+pSuZ
p36mykAUE/qlysXB168Iu9lvvcu1UzPkaMLyBvAJe017QnTCoXALb7In4kmen5Mv
MMXGj4Pws+rN6SKWTYzydk83GLbRdbFliYKf1i38w4vNKZPd5EwG/gu7QF5mSYK9
f3iJoal1xxJIih/wpinkNbAWuGM8iYo2hBaoYdoDlnClNPamPG9cUUcME0iK4Tx4
WJD907lS7GscWGAHP+lBPW20ye5pEUy06gg+lp5FzXK/5LyoWEOz/MQ3urVM1ywU
ayK9XWjQVap0rDsWcKs0vhdc/EJFQqEAZZmdf46J8jXxNaD27HZcerzpwbMrQ6wi
q5YMnNbHB+0pZDFAoVp9etAu+JB6EdGIB8yhbUUVWM0EOcaroCbr+YfhdJVdWYKN
to3L28hEJgnO+fN0QQQnRI6FLxU+c6VeXu7VRDrXOurcWIJnBH+hlojKZJzQ6fOf
Hu3n8vdYAgqVFN3aa07hQ2ck1I1JsVZshgF2fHvRmkPKVAcPdpUdK70ItFg+AOxv
XNcsSB2llQxu7m/K6VN8lwOBpeJNhi5/ZnBqYBCe/KhHd1sEBU1SlG5S8uSP/Lgs
r4b1xP3XtiYHbRS4j2Pg+ewO7Q8xCEWSXBlFo8PeqwFQo/FLd9ziuFDBulvz3Xai
5MTHi6wPOVnN2GiAK4v82tSAnZnttc62FPbMO8gSfP0Oal03JtYoKFLxrhnC7T3w
b/tSxh0YZxdX1AErnVgWzMGdQmvG7P33bt8KQWG5tmz0m+lTzlikLmyPJsG80kXP
4X7da8zPHtMgFb2hAysOSGpkHT2O32Ay3SsarB+Aix3XFGJ1ekSOyGnOtN9Jd0zi
JeEG0E5zPbpUOaVl/qFxAurMgFzqtChcfljWrTGLBODZKBSKu9ZCTTuGgK/Ix4oS
LDWaPmO1WLk+uHYRp5PLs/s00wFJx4FpfwUAoqAGRoc5dpTXVZ0MH0C2BcRdfNpc
LnbptStWKpWyU7WHDN5aUtQl/xt+CsSLILXGKLA3ON2P0ZJmmdTLlQJpWK5tCMaC
lZx9nvZYkPMDymHJ8l75ARkfr1dJaNtMo7GGNfA24sd/msbcWWY0KFWTsfEOPXEW
upw7/1g+q5X09KjPNT3ktt6eD1pYAR5rrVxOnRGNGKk68sgbmtzJXnPq8vj67r6b
QLv1qGG0FTE1V0HxgCCkwGmQbJzqxZgG8hc1QA5dltIPsTL9b4lySgtqW8RZFEFe
k1iRtO5TT6x/K5OqBoh/+qvAfF+M07OMNSJnMIiIIfMCavGBCp/UGW6OXsulm2ry
+m+eqfkJzA0FPwq7hYD3EWAGkQZd/0+wnIXPaR1/qwrHT+sEjk9m2Ro+ZnqNInQL
azRQsgeHhdhrSkodplK/6+tqFqDbY8jvzIlVAj7IdnYZ0lB/8hUQjlRNcDJ51Q18
7IPmOyaO/aqY5AXs7ILCuocrZcsSBneUP7kbf+KfRHqz1lwesYQX5KLBt9GAz10Q
eU2wgabKP0w4k0zEIiUfrmTczglbQUbMxpalCetl/olfEJ3RepC50kdSXM1oCW+U
rlj4cRABt6t+LHMfXUS0lzkLB5Nb5et+6q48GQZC4LhK+WwxVacFWuCUsUSWLj2Y
tj4abILksDuUzYPES09pJTjbxJx/i39EAqD/G2mk6U6M3utEYPbpbNT8oSGQJXX+
zdKP6KQuyQiT2EVHQN2VCMDQUsh5+ZdRPzuXksUoMI6ocjPrZ9nSFAnBS86wNBGc
tWMYaBUmDj0ThmhdVHphaBRjuJaLNnJ+2uUQ3R2uD93DolgOt3XimEjDA4W12V9y
2et55JTT3v9rF+SMpXDoOk+0+8lonnvF5Nio4ZXUiyNY+M7aa2SASYJIZzGh76lG
MxRGnzetp/smOsQXtJnCYz3IO3pqqfBCsYS1IeZduvCOHR38790MaiBjwFoCcGD4
TiSEUM9pVkHeTnAU+KkeFnw7KBrOzE1oL3NtAlz/262fiBEQHibKVO53cT9BabwJ
HJo8oxq0+lXNv8ijH9WkfER0ag1EA5orHTW5V5KRB2aKau5CZrAYR/CBqL8wVBLv
3TxfQaiU5+Zd/HPT8qETpY3Vkd3KnvYCUkqRNTQ2HEGHyzQDxTlUgz4U9G/eC2EU
35Nf7O2OxxdkbVfE8bMOWrS07xQJaURuyACJxA3OpuZIiI/07x56pSkPzYut/vUp
ZHkGIQklA4iOgj6RlxgFcm1jaDUKXP+eQkYri4fTqbLy+LJYe7VYE1GnjL4Q8xDW
XvXlNm1IQbeIuiL7gr5WJX1Ja8jSasRr3FRuQqzpue1PMMrl8uhn1T4va1l5b5Uc
P2RjbBGrzU3PGnOcvuCtkc6Nl6ormFfWoBY+llwyM6mb5cJZdzDyh0uQslPdL9U+
SYqMp1Q0BloQuwxtUSmi0eByu/6nt2xyETd5jCikd8rnbnuOCm4NiWIg745SAJb5
gP3oZX1QxG48GrkhJDE58AJe+Z9KJklvuXQb05KFK31AYTrD9y0xf4gQM5wPaaXY
YvgK6U6i933Qw14NmH12IeA+bU+YkSbfPi4DygvZbOlqnobNLpHPWQLzEP3JbjBd
zZUwm6jehyWoerUI59PmOnEkwwNsnCyuru5beK6AYth62gNBcIsbk4SgmDYktItx
s5oj5MSTP92nyHytuuLdjrM3UE9/d0XkJ12/TD7R277DVxBlZXlZ3FUOUM9LK6W6
rPdxHy6JM9xGgI9qqNeOvKfQCx10W8i7uC1BK/CISaG9RYC5MmdCG6fcxXp8kMCq
sNHknVxz6hu+cK1vDe5HvbqvsdD8SwypkGQxLLePK/EhMbjHM34qs0uxdwmy08qf
zpuczwzHa6jnp2MmFVT6eSkxsX6B6fNHV4kmKlnCcgSptgvP2b89cBYu3atX0Mh+
amkt2APxR3xmM1d1yuMrOWKaOuomlpeFzNXllwr9pj+nR8LvZgz3ollOQDsSRQr9
cQTYUD+IFw5lj90Xgy535Grm1YzAA54+dbHk0zqA646WgKRokY30tVIsU4IpOItE
NgepGz3Q3wP+tK+PQYrd9EtV5RgtysUzHZPAqTdk05162fAGPkKFbvH3hh/8KCb1
Qy3uyhnEg3OecI/54srgbAr1cOshE8gi+//sF0VDQRE0+zn2Kokx8g+6PgBBhqhO
QguPBFIg8xJzuAw6b1zpdFz/UKmItQCmft+fUtJolhD+dltf0JANVviS+pNIpWOD
khsznRBBhhb+QXTjBmZkWBYDTQixZ4YP8OyElgpepHhR68ArjhHq4uZvTPfIDM8k
d+wLjuxsppUzZdxN6fPAzobwllt0u/bFgCuU6VbDS1QHVLte9hmhp0+cxZF1ufIT
hNB5Ql6W2BGB3uwxa2ScbGMiNT2HuBlJ6+3Zd/lp3VJBxVg7pZsncwNss2xk2zuL
O7fOJniPHUaZJ6yWmfrT4Ut/EGK48t594XZnfdEUWZXIOPwY4lkKRIgSzRuUWuYI
E10iuuN/QpgBk2aC3K7PgwRauqOcY/ku5XYvxjGCOj/Tx3uuGXQoMRKxSdus16FF
BTmlp6bsVDnur9cr2lTaQWzUFulmo7ia7Nb5i8UJ9h3OLmXYlt7IR42DM8/qYlgd
AgC4CS3M/AsdJHoS+zgC2GQ5oq0quKJTczTKA8v3ZNe7Ehc+vPCD+mT/kcfy4HJS
ti1LkJDX6JQiuAaOO5yRQIxrKJEb0TcIKv8/QrBd0vb0gGdfkCKM+evQylDzWGiY
PosR/zixz5W+4mpiV6I2FgOWX+vKnv0pQ0eTmlGn5tdCfIGGLtzcboWeT4clXlPB
jX/Q7N/pqMnjzOGJbJp5r7yzXfI1t7DpSkARv4bYPZ9Rv70Fs2W7L+7h3tu7gky3
CNNTY7clk7dZn8+H64HRZ3E7bN2qVVYLhjE8Gd9WgEGY2J72IUZ+4uZm/NoEZx7w
lq4vGX/63SMwzDfjnvq+dgNlGgCjz6E0Q5KsqKzB0gYw1ZEsiZV9180sISLoOa6a
++M358QsiaQiIqLVnjrrNtpG0N9PZvwmaR1aMCOOplZ2mH1qAXiegnHs/JsJfz8x
uOo6Lwzu5dky9Uo54t2EF4p5jwIi6/h1VNLD9AWZ4JCx7zKfn9QE5KGX9exuc8dw
7z8PYDqb7lrqsuUFFoPsYZkL4T8qx4OkpgYwSyh0/ykECw5E20feqRLmzvsrL851
WjrZec+DvED51dlmyLo6wFa+WB9nL9ARu+J8Zik3X1jnlnhsgg85yRRQavDQyRfs
98z/GzK+QlTcinISylBH76ibnepZjjpDBAfN8mtcNzM2hybbFs+RSiTkiKjM3+DR
HxBTjuZ6adb8YGtQvkhOUstNolTu7HaetORqCNlV6eP2HWtgg3UukFJRBHBjkMDd
4d/eR+TzMLxSNRDO2cr4Gm4nKT23m/nh9HZDFn3UcBjYB8pgv+ceMSX//q9ERBy/
pVvyGQRUDKI0X3HHvnOoNtKCSC+epWeK+0/FxDn2n2IcMQ/CViUE+NgO9k8ygNzQ
WhOzfNyjOTCi8NHV/aFxVrTpNeSS9nhk6Ywqw880PGf1kQgGcCPY5PHkDE+2rIVy
z5B5sV3SrV8LPmQ5UFWmp5yAKu71B1v0F+sTnUpXwuznXpWoBczwkQRKw/IEkwnp
91RsiHvxGfjpOJlvdFc1iKTem+WmEbX4QGnV+p+3xfXpU78958jfb/318J/RUXIY
TjYXbw6/oBZfgmDB78vOejwGqEP5dQNuGZ9DCwTze5UT2YLWq0iX0gTz5iX/x1Fh
dNf6PnvsZH5UBSWam0cH+LevBpF2ly95U3WTKqrJgaeO6St3iwfQlzjB75TDA+uF
m+wsUfbMal5NIYnxNs5TpmEyszOa8IBC5vzLq8bARug/GZg/dQzM77Dwb3GmS1+E
t2wGxbvIfPmBH9iIEFOfUacgnUS5mbQCS5IgYhu6cDmTC8TR+t8qmGbrWN+4j9gl
NrXycqajtGXLTIJDi7b9wORIzFG6SHaye9Oo3VVLn2I7/rNdyOBT5LAcOtTZ6wMd
X9N+eC5PlyjsFvaUSQT7hN5J0tXJfbOOnS2jc1D+XdR78plFaOJFiQr+c6DzkxRN
vvCw+vY1sXT4UnWsAI8EBMvHPJQT0nR0Zai5gyc76smESCqvSk7QluzrQzuDytDq
4XkeLFlmDg9iL+eph4AgeenWpS0K6w9Rp6CtJYkAK1gphk0UNLD/OWxywOce8meX
1qwFdaM0NICZwaL72wKTHgV4HakWi7klF0CXoG/SlK1O5cUesJZ4qd9/Qt75dQzC
AgUJoq0mVistDQSSKgP8AsYg9vgDeEPlAlpzAxPU9qFUO9dwmAe2l679QtvI+WVP
r/4nQzleW+w04OvY/t6exTAk8PhN/fi3zT2JwMvT+VH7NbLp/+Ygj1ZXX7bm20o0
fVj0X1VJaknOv82nxbN1dDWfpt48vXMmjWShH82Ame0JQX+un0EkWzZ08+piTKTT
zxdhhLeqYqCuWrqUfRNw7qqEniEAytWou07EJtfUJL0eg+8/kmB9rcJFZqdHLmgX
hgSKBUv3CTaflPFGTrwjmHyDO8hkf0oCWY/INcCI14n67u80iCUmKjpfN7PRvHTh
EGrnTUKjB34bkMm/FtHzNZUjlx+OVnyT29x+SrJRdFTB5evcM4sCVlbtmNb0x8S+
Lm6lIgbFR0u0VDTJPbsij1p+VNrf96tgFJ1iBXFhLj8pidHUPgmy845Z94JdnvFH
8dajc1sh8aIdC5cKlSr8K9JzDa9lWQ7mlMSNV86PbB8+rZmuwXau12Dlg0mMuQPH
RSIr3IzewdTDI4WeZD2OqC/eDCZBgrmJOcyNnNB7J3rcBw7k1NHw0ZPkpWGFDQGq
htS3ey+yWtZ7xWoovKHcRFY+ZuH96clTGphyM8My2vHD1gvLJvwRhzRcQrAf4VUF
mGRiBMBXQxDtP9l2jdjVtcf/LEmCJupmxFJgA6D2DL5x5FQ2irtIx8aFrT6ZSB0a
2GrENynF0SG04HnugIIvA2WVNFFR0Hr/xByAILVKJmn5RPnOoIKrWwnP35itqawI
c9z/8RWbgAi0UdyGPnOPWOSA5WCd4xKsHsA4xicAO4L5+CnfC9p0xjsKYwPOECcI
Gl+jkPpiCQr014nO9Y7QSzIN4KpjqMXxHO6CVwGGjBNpayYO0Jr7E5MPP//SenBH
YLvj9gvSp4Ba0gyHV2Gp/CD/yF1DUE7kVysh1iM7exCa5f/0zNlat04FsWP36tD/
3h4JKL6Q3BpOlYUQJiTWiN5uYTvjSi0bTO/asa0o9wVODDOnr+MVkhRQlPOfSsYt
5UI169+qzRRKlLNU667hBUGCSEYLS5dz96TJqkfTQ7gzm2b2FKDeIDFI/hF4MPvF
GYEa39hufS/b0+QTD21RFCna8tUtmAjeTnEhZ5e9RkZ9IHieYdJfY3uAsk2pnQjN
ITp4xzm2wTVHCd+Kr2vutUn7qbN5vUP2t7ZP5uPuhZuKRpGkwe8iBqEJDFLYzYza
sz6UAF/KyafIcX/mJWkm68E0t/PE6mlOSGRAPBcCqBM/AHHKZXteDh27p0adXFel
Lm95Jyt9y5pOi75lf/vr3EdwBwjLh/oG39d0yYlhlWr3Z5jyzplip4L86q/5EpT7
7/aoDyulfBbqWGkNP5JstJLfNDtlUZC5FfLcjs3MZGs6hbPm7VZK4yYoHdY9VXHZ
QFXyU659T1rIxWXj5UDGj5ac4Zivgggj3ERyM/bhm2wyxlLQWx89cYqKApOabJNV
chK6VvLAqeqTUcZShr2R+f7oE0YdRuU7qbOX5ZqdxSYETYTzjCLXchzYD5azeJc6
HkGGbhJWKgHgL41L/kMinKNJFHXIf3GVzIfKmqKw/M/IAJZyeZHTH9TMyYz+Yhck
PN5XFzdEOqrFJRRZ4Naj1GhSGFD77hzxMMO/kmS3d0YgoJ2LsJkLoOFUvHwurnHH
3C6aO4rJb7sEkJhBjuKbG2E92tY6As75tYqW/f7LohycVmLI2yWZBVdx+8SjKFLb
/hZdUDlsoawv7GQxLTJNjADHpUifNrY9VUZ7rx8S3+giEAGTae/w1R12GcXhncam
+OoO3psRsFPY2RzXsM6UU5dMGkT+KBrnrwCLx3J440QHuu8S69XSY2S3HLhrmKeE
2xbuOO+6lJ+CizPgCB8kBjOSOsJtIY9XdNgQJYOG8Y1V0xsKr1AwJHXxbhlrFfS5
CpKc3HDMiJV7oFUWZTiT6DZ7fE8uSKcfyRHhWLMkcsi2i5itv/yX0v/S+QN47e1V
ebrhhtCTMCGGHgV2MySSrz7sVsQ1BC68n2byiE3y4Vb82x4nhBBkowgsw/O3id16
9he7fUoK5w2PmDjUH3ozesQ9WHod1Q4ZdUTfXxno3/mwHapwPk+RZvT+yc+vsKEe
iJ12a6NjtImqcj9YeX0eF/jpaUc8M6KTgzu0X2S27FVcicW9UVUa2jW9EqTug+qz
Siv7pU8aAIyEF3pg1ukLagWcJDKcHa9XApWIhplbcm6hzXuaKjMeRXZ1l6wSA2JO
WeRjzdwJeRXXjWZ0q37c4nCxq3rfx0dGW/y+Sv/LPZ3t+qdXL3mVrlAzWCsD1gVX
suvk25qGwODQibekQwJ7jyD9aVssg5SdLWFpOgxrF52ymHNYKRvXDTYKc5hTMUCB
G1k3Q1DfE9FGaLJcfsRBPU3mKtf0mM+00YXjwPhuKWZqsCRkw+NX9VRWJj6vvYO0
FiT2snozTYK4eVvpX75Ix03x8Z0iHn8CbWD8c2rRd0KL7u8Bf6PwVrZb4KTNNPAq
3GftCwn0/YdLjEbBiCajqOEItc/HNPlkpaI0eLkPhheJiq9FyuTT2BrJfH1d+OXo
CPs9rZNVAglEAEW080lRPjk2FphcDzMGCoqt2GenNRCcX0cOsz9v9lRYRB2Jkd9P
WphFMPzWYKx3lVEy2hVJLYwA7KIQzJm8gOmDLB8crfxnldCr6eTGozpve+og7PZX
jvjNMn1L+buzAet6qD1wUMbHpFwWrcQUAb9eRNmUsnkFMJHCbftyMfGO46Fw+YY8
aJyTI4RV5HtVeog/TmV/jocUKXy8+7C3/rOCtB7FstWVUZe61F4m87QOPmSvGNZP
7ywzel+y8RLUy3xFDvPK5HBR6d1fX+GdjVKPAWVBmj48t5zgRKQoQ174V5FdYFAZ
Zt6Q1f10BtAEbfsdYzqoOQ7kUk5dX/eCKjC+Yo38n780Pz45ZzEvNSyYAIa/9xXh
AM5nAqqfdGVVxjNzxytn+uNmGwejTUzfaqQBzF4r98o0z8etStuBPcmhsV8CPndW
vKQla4l59uyc26YzNDWbsFh9BCXBGNZNhaqEeY+UWc+P0JuJmtcs/RFBlzftNt9E
9787aMW4EUNuuYppRQnxcCYCLaRVyOcyhl4ZUdadsM69X/T+sBTDRS2GfW3wNKV7
ZO1ZvDAF+v6xkdb8Bgz/fPQoT/9Xp3IbA1oLCUonJRm8fi7HcUjOkHTaWk6kZJln
ck4V2cdEXt5BEhzaJucNiXJ/BWF+IKKKuHp4AcakpCiqXNO4SmuKg3DwADu9P8MV
eMUDGqjvwkb8m8+t+11+Y8FmvOlLBT1HeRGdg1gB373UKtFL1ik0FVDzL0/u2wkX
wUx5LTcLIt7U1N8bfB1F6A/OAuxV18shb3KrfnlmiY22k/O9prUBBbX05uAxwvYK
Gs/IrKg+DXipoMCiqB8h2ZoSxV4D1Cfz4YMkfMwGYG24miF36LUjV5eklsbmEcf1
czDiMdh3p7dIbOGuju9LeUKngH+jn5TfA5EQzX7KxAfRH9LCfsEAMwwX3mhNAPR4
gtHVTRGBz0yILti42IoGD6xRVBBbOcbYrs6JWMt5kV2KIWcpr14L5E3Snhm0QZZy
nRlFi9RPv0jTrgBaegpwFKcUeByWzW/PKBKnduCK4iupa3mWUMEaNNCse+8KQkzF
1WW9tP0vG/mjMeHnrpdEgRO/lo43WjdtQYSjwPbLhOHXjuZMKVtTNxh7JLhLlfnY
8tsMdv5SjHJ07PErHvL09xmhp1N1VN6VqDuECOnJYM63dtFu+cB60GMeLS7BE+gT
VYYeZ3l2pxW6wrx7lnOAXqlUv2G+4aOybGOL8T0i572u8ZHMmIMIps6QmD5K+QvB
u/D7vb4UPyr5bezmCwHWGpf9GZgg2nkgdy/0kmsoWbMtoKVvJWG9Pmss3LwCYZC2
ZTKShWlsHSf9Q93JB/xonGoltmdBZTL9qNFMtzyF/iXHelQOfSf/diMHZ9P6EqET
R+UGOXVjDXOpvxZ5wk+d/cpQZEkijPgZkjARetsfcDm+1f0rbmrnX2wucCffU18C
dAS/mQJnIeZyr2pyBKXllgyFQJedFg4KzktlPWqVhZoMX9++bRuSFX+n/SZ8y4UO
zbHchpnh+bszQ5gAh67rodggkTfH6g+KRgBuCxfHSINOPtwV6sM+ABoLKixM3Tp1
Cc7TT6NONYCy9aTYxVVZH3dOcvfFsWC7UMq/So8dlsmDZVBuLlVsK8lQi6Vg88yW
FFzxCIg4Adz5J5+/YpdMfhVWP5HL7km5YzUO8jsPBuJCizhZmEpKlRLmzjyL9YB9
mhz5+moFVZLkUZWCc2hIVkw3ghtSgwoHGGMJiG8drMznr3WcQ0zwvJJyQ+ppRVGS
lt5TyrGwdZdZIIsimyeXju3tBc1p02jMTDQT6DygDJl+ZHJMnyG+BlhE7agBVp8j
OS01lse1KSb0inNM+1JNk/9SnE63ZGWXA+ULOYntsZL/qQFHI9L+1X7+30SKnvVW
p4XjalN4lXTjVS2AxY9w5RdzmrSNTBlZAXHp9qSPJ93InKbQS3EkD1SuzdMhf2mc
MAv0RJCTA+Djl/PNhiHGvVIP0/AMoeyX7g4YXGnNp0xuIy4/Qlz9GxArDlSDe44M
uZ4OitKcr4p4ukpWZSPyWfbt7oVdU+stDn/zvLLAea1wCDPOU6Ew7I6PHeB6sGKp
RH3Vq+CxivaSecIMwHcVYouW7zd3+Nnb1F8Fba/HzE0LkBz1Z1hYVQQ0S3pXimTF
YdsNKh9WO4hZ+TwRDWEILWqg8pDFe9tAG1F1ontbAScqzpicTyhjGY+QREO6Cno1
xe+DjCqPNh/2RKwxGq3A/FXJLJF3cHWGnJZHVfw2k14zDkNjt7pi7SOVQ1lrwdGS
ZywzfBnVaKjD+iyKirgYm9XifseDIotUAPigFbtiCkgFtSBZ2BxFGHEAQXjtppZh
Zqc8Yp0s2Fe/JauxQJz8wg7m7yhT8vn7wxkL/a8/ZQKFJb92XkJP5hzy0XgI/5D1
dGqp3FUouua6iItpZRDGZPoX9vvgTM7f7lv0oKwLjx6CXhhpLqZwM8qQSN/AnwTN
dc/fN5wHK5KEf9CKzOSvwvsnKX2J+PeMzfZnD4Su1WZF750kMsvwg3xSkkKflhnX
J5a/Y6I/1vAYvOwwMT+M9yGMSLCpsfBq2g6lYs1iamph/j+N24XFowc1TCWIvnsE
5JSnrw9dEAmpvUWAk661AKsCzKwcZ5FOPxzMH/zhBpxPgixOTzCgbmrlGfq0myZd
3zehKti1Bt0LpxlJRyI6TYh3YipCIFRMpfXXPKG/eAeuINTLiJpakxRi1YVW/JFH
wIYJbDC67QWBkoHtNt0tCEylsm0DJxFZeWjY5CvjtCecGGvsRvz8Ex7T5cGk7U9q
eV6jR3TwYRFHmazHmYg43nW7z2tN4XCXzJNdqSejzwfsS8KA+UWdV7Z+qBSxt9Hw
/PwA3RH+uyRVuIctykAaf0qSUmMGz3H/r0nkoox7d9XfkfqpbXz2V2SXIpwTUnSJ
X33hB1FcDie2qBCYleeODUb1OBD87/IvofwewsSAI88EIUYKu/YN/c9G5wRcm7PW
bOZ9MH8e5kwyDKK9q67qNI7R+zOcOewmgwXN0A23miFkCChtVkaONnMSqV1YEo6+
dFhW/k+2I1PdqjNnJO5vKJg5IPDoc8x4PChJwvNc/yqVAdiBi+yhO07DM7qfzRu8
Iqo7UM2xqI8RtvWZ/828ByQCZDS7TPEvPkeILmBZLqfyVcHQ6kGg0Pv5V1OqoOwf
JpVhrcy8iAUJvTDQgx5015gloE3nB+fdSJdFcbZ5uR1QCOsqiK+R77zfamM/cAJz
2jUwmZYzG5s0SsffmTyNcwwUqy2TxniK8HGHD6kr/7PZKVl0Ykl6l2sM2RRi3VtI
RSz+S64bVcqvK0TCYeZUdG26K91Ek44aOWs3k+29oKYI6Szo1sX3T/0I9RShE05x
sKweE9pzR1E3JrNSy6FuVRLaZt5Oz2XHQYkcLIqcRrIrLrH0+vTOny+4qMegzgR0
+RSX6ZOhgutvSDEZAScD0ojlYVSDljb28DJE38G2A0a4UEYOAeEbKafJ0IOx7cIk
pWFcj1k2Cnsj7OdFQWmQW1gqTwbcrcQd7xMJtpVQp/5TFu59vfNQqiJAlvZimbVN
G+hstzqxudkeqtX7SUOrbCB0T3C4FNHiWFD9dOoPhIPg3kvI12GbPXMRP0c6/Qht
TLT9pQiMzqUPeWVylLa55d799R8dyTcVKyjHo98C1JPhfmY4zGH79n/ASuy6DlOo
BE9qj43iMp4+hQNjaCJOKdFx3TPAaxqQnvf4bN5tgresh6BqNhVZGcKMDlRzib+3
a4MT63Zl9hk9/ldhiADOCqe+iuh8lb4H3KSWzRtRPxWY2/BtIsyx8KszyjGhMFz1
hwo7psS41r21ZLGBtLQrovenNLU4EGeOFbT2liGz3RaJAsn51rWEkt8bLU9dPdCH
CcYKm02LWDCsLd6yo8fXwRCF4vYS6vQ2SczjJLFfNDfCphdOEE1Tdy2OhqGxv9Ut
CJPBQP2uazhEkL0soO2nuvoFwyiW2V6ZoYnKDeCfVrOSA4YjN99nNM15yKvnQ61Z
zz3IZNMK69ojJ6OcjKIZc6f5arokj0ihEEIoyOto/U3BSvJb0PK66VUzGWO2Iysw
bFVZlhhuwcezQQe0u01vAfCY0fFxmW/gqOlV9Jkd126LWRT+cqhhr4gi3SKDDmfM
n4VNiGcPNTB1oG6FbAm9Eqfp4/ofUvmNvQLK28En9B8bTVDsAKNCBRG7UfqhVvTO
1K88tn+3rG4zgQqr61GknAwtdezW2O0QIZe51msaaG7/hBQVgm718cREQgIq8YDE
gP7Xs+slnyGAJdqjb4SQvR8uZzVt3xXLmdeoiTpL754GWBsGJtBf6vRwOS229LHv
5RC7OCtIHb/y3wooR025SMMRkrzexaN8GL9i0fE0e14DvOdNClmyCzDP9LYQu+Z4
hjUQTTXs6o+qfBDZPIdh6SNZDZttWCDR8tWnqFPFIHanh5W1aHIzAvecYyqu89Si
8NwTaDjHGkvLA9DQUxc3cTIfuE28dIQppSVLAsSwQWE0DS5SbPdMmkq/hdq/+kUP
jTjfn+3zdyBgdVsVXZ0YPKgEbtxoWqXm8HdIBoEKo3MgmHdjg+9jthfnHdRc8e/B
kggOQtT0VXEC7lMuUtRgKlG5NopXJccUVvsp7sqNitm0EDwdgkZSSfaULMPsp+mC
Z+kx3AqTPGWb9dVEHyE4G/N8QXd2+JQ4UCLvS5KApeTgY9c+LIj1WoH5pv+nBri0
Vys4hrA03BFO58W5OQ7rXXAaDCc+I2XEt5OvenvHkmFnjtBVv0m3tjhwsYpDf9cP
1wLHoc+isykOBDwfm6CWlCsia2fmWgNVYJZDo32asEEM/pvUGMa9ezLhNGJaLrh2
bUvZWn8yNyJ24wGOwUozdAd23lTOdoV8rNMFzmge5hK2YB6INaObD75kOw27yfH2
ClQF2Fsdoq5f8rerkg9Xru7+2CkZFJoWd2C4YQ5U2oeVOBompIIL8KtUdssmFtzd
WYWmhW5w2NNSS4IMqt+FldSoXX2aVrEW8HXps4ZIuYPMjCEBqOntlBz3R5z0cnyc
QenF+9bYNO7p6n2nS0uw877UFiJQtSuSkSZu2IHoKT199nWQLSb2w9YnPCwnbDzo
idBrH9JMRgU6KJ10GgmuBdXXivNFZ0JRo/5wN/xKTdQY6iMvcfnEzdFi3u9HktTW
xm970Vv4iiEu0axuUcbzU71kw/bAAhWKBc1ZmCtotg0sZDSVQSg0FDu5liHXu/nq
nl8BdRXIKazEe8Vravzi68/noccVcdOOE5isFkSAZaPkqPoJpoamb6pQfjSG/HY2
REEGS1QCPrUJn4+UIONIW9XNLwpXRpyaFqCDNMR48pYKA3dXfvhmIxRaOh13RmBr
NLj1K6T63nkzZLTfL1PYrNIs5Z0cfRLhOV2/jvck1EeuvJs2LaBlzHTv10KA0W+Q
o0wL6m+bM6TrkDwiBSpqcz5awUB6JmAlfGgnjEHXCsWqt1MIgRFcYd02dmhwB6e4
dc9Zvj11YWt2oBDixBqLRtxLj/mqQFf1B9Xr1tNP61VIN4dFZfB57hvUWvYn4Jcs
L1tI3ky0ghPC5BrWrCORUX4el1DqX3/3ag50jRiTUjOOLt69oVCF9ghO874rsX/q
qjEVdmVZSm7YjDLWDxsnAlM5YXwI6WOxZxUBo+CKDwaM+q+DYbG+zBl2mr6z9FOo
mlEOAA2N1HQRqD6l5SlKvSmdbtjBlgzwdWpbVv6mbCqLGO4Js2pXq+CagUeAGblm
5GRYZybirlXhv6i0yZwRmT2SzEdCRq05wyaRj6JapTl39vli+JS1GDF/HGx2BLFH
fF8xFCyi+nFWYVQv2g4Pn1gDnbj2G9vhgLiNKBoweNMs2R1+WwdyTJOnhwUtKGgY
4CqH0VZ7WNZipsA7HkEMB5ZYwC+0i4n38h3HzW5CkdHfrGnZDdo9tCOhEMX0mHDE
fM0QiAEmk8fv71TmgP+mppATnH82Tp/YH7O17j/Q2SNGVTdcpXyvl2O1mvcOpii0
fKmRdLXFuHukX8yGV5VM82QM2+UnmgnfIh7BUv9oTQHobDSw7eET9kTydCLnLvtX
5bJP7Anam5VqMLBwm55Vo7+iQk4zkryBfoPPhPT3xdm/CN27arQboKlVa7CrT7Vy
UoCIXZhLZzT94xrTdGb4bdTr1MQyPJMU9FZZEkINXyhIUFSOCrQikMF0OcfaD0+P
bMBuV2GxmwZbpY+wvHfJiaXU9nXFDhu/ng++uqJgUJfjP6iFgMMQoxkMC2BBpqKd
drND6oDsVGvNJEigyruwGv1rQXlTm5pknulDecR0fRgOisan0LglkG4F8DwJMCA4
boMZmp0zvpisrIykKm2HORppWYFEY0G4uDhH5YrEYoLVcmW1EIwBBsiNnFZe4IgW
ZlU9/jxDVi3ODCD8f84DC+LyoD69M4MO8T7nRY8U8qo9L3+TBjEb72o5SLb4cEIi
jrbmjzAXABsyg3iF6VChxYBmTF5BWXAjCAvhKFVj+iFSbxayFaQN+EA0LKCf4hGj
E2b0pPonN0iNVbckCeAOLdeL88j4Pw73Htl5g3lPI3qQr1TiQ8KvoOpiqScM0xCc
lE8a5dwefnW4HCJuePYMTSK+aBShV+bWCs+79hDJ6oR8xGvTUUOPEmFnGKyqdVGK
9bqeD2FPkuvzkprvVdsfY3hmP/jkGTCiQ25ij7OOKTmsmI+eIsSFw/HwBaSgrkgt
ekAEX3zzxqnucql8EW4JHLgCLf9ElY4EzuV/C6S2b7RZezCMOmbP7aZ4fY9k8bCK
mm4VulyfkfksIbOveJSZ9QiI9T5gIFak/edt5hdJfAxRqrvj9rViitSSCASHMoO+
0xAS6Vk1PewnjNfeRhhoDXuWFpwXvVoDqrUCK5Gyac9PJdFM26epFKSyKPtxQ66/
jGbMaAu0+I0pIkbC01Hr8hVaSXISuMjIobLirCOYsE3hST2s79XzY8xjuUAo8A00
j4iz1ng58gw4OGt/8t1BTKe8FXqXT4Om5xagyuJEXmykqNq5gojZo6/AP1O5di3B
KbJXqNsljHIjsTTfi2Z/txPTwX9W6m3ddDec0H7pY8I74syu2VvK/GlEUm32HNzY
IaXdQSHtV5OgthVuV58vEFPLTm7ZcrQ0A+ZFcTlPL5640aDB64elc5BwnXckMpTa
YGHtsxUCusE0xzd8MJVtji1Wc3ritahP1cnuUCQj03OuhN0JHTWgPtjnDi3w/4bA
zPH7i24lrtinup0uoGdI0Rq0FkyRrtq2lP6dReHvDockgeKuQAz1SH+3+9sCu2jQ
7gLe76WTt6+Peqk9khy3msqMKBRMMI2XABjSGBmkuPrTyT0kEOI9+xkvDGXwTr0U
k7U0I0D7jkX40/2KmgSAva0lwPA+pRxHwL/Kg3l4wq4Ni0fFGkw6COoTh2l7ujmN
vReD0s3Efir3I6COnQT8PnBa+hLCqNtK7jST5wTbM8AG0MLuGo9JflLorWI/BYHU
49Pn7b7imWghLkNnAZ7eCHBrjaTYxS0waslOFfjMeXkRp9CJc2a9CwP0ZFE5g39n
1PSi9MbtJulJ8kVs8031Qy/6s26sWU6WvfRtskgowvDgn+7GhRpyqekkIrxITIEv
4GwpVNAVirDD0n9XRSEpDbrTYTnV1zMvdCIQH8DZCbnOG3NnFplji7okzFAhmZ4R
in7p8HBGgBTjWgNRIOsgbB5COTAcmctC6HBUbwKSIJN2IoNRO58y5OyRqfjop4kE
u8+tYI0vu1a/xrLBtn+4+CRjxmbYJhc4gv11ckqg83Uqq6qleZTq5P/9oXJaEGoD
Dn5PxOUVHR6n04yhPLmIjZRnntcDxzU7OWoVIvx2DnqaA4FK7yGyusgPpQK9JtgG
BGEdVfLXJKKRMH72s2e2fmtV4hlwpC7166gSKl2fflrx6m5m/PfdIoYnEyJoixr9
/vZDh0QJFKvFfbtqnw+QNi+/b/D+7iycoJLmmfUBQOTEac3S+A7gFAgDfwCYTrqP
uSOvaonZCHOTHFfvcdC5qS+Trid+tmrptpZwbslIpjTn2atRd4Shc9hA6ZTxqS6q
gy1gWNNQJUlzv731XGgEQLhaqwBFgVZE44krOG9/TjnN9OtL21rs+FTCMbEHEMCP
CRvgm8HDezVgIeTy4H7ddm/hOCboejsClbF+5LZs0LS9B9+FW3KWQ85/A4yYOniz
k18C5T5Uufy4fK0RFWdjZI8lJz+EfTYkJT/CTO77ls7l+m9sBdTlfQfc1EFTWj07
OV3/Xn+0Yyd/dgdQ20GA2lRAwLzNsgUpcjur25Cq1jayk7JAJPVa5KjxbQLuXT+V
k9GvQCWzFEbZWzaqqfX5OvrNU/NSh1b9KOFN+q91GuSVilySOdJGLTcUtr1RZeAf
lK3MAGz3V0f3LRzJZTpbUOaTQJjcCZbJl1xKTb4V2JC0BlfNKx8PjMxO2cs3W8L6
L1nxdQBfM/KToapMYc9ydb/vMK82JYzl1e97NtNpIko8noUYv3paMsxBcHniKryh
jPoClHDQBZxLYzsvbk+yDohCW3DrANj/LsJqIB0vMVNfYBm5ltYfhLRLgwIaByFC
eNcmlGsGFfRkNkjFYwcCy33el5j+z773tWHWXBWPkMM1wgVMt8ilzJGo20UeQTR+
2oe9TxbHjH4/MNQAXiI3flVwkcmXHs6vSuEfWoUE8YsqJ6X4+DZjyOAJS9sp7ksK
007qjB3EVX95ckVE3WV/iz+dlfnfu0hi8/RyoHfkoeQbjn4dMPSKeDXBAKUS2uDr
xGCeYbtORxePmuJjnCRwhD7iIxWuEYFrqFWnwT/67BI3C3pJR1xDkhjKcwsJ2uam
RRlxIUzEOByGCpvizZjEsUN2U1pZvDSmGaaCBl+2EO2PhMK/0WEqq8D+3f04kSD1
SmP3RM701Poo9PvWKKAxegypIvYMe6FgR9lFwko8QrMdUa6EOe3Yy7KIpFJYbQKp
H+CfPZ4DsFczjPszEysQ3fGad1j85YbRP/YhmqYhsZxlCMtwEdcJ5a3SRE5WF95+
bgirqCQUrBpROWgty5LsvrCqCVDz4NXMwKgkgeUhU1/45dzo/kSFfSKvtcbfk3oF
z/XLL0DxxeKXOw5ftInz1fabTHtVB936sCYMus+UHJPnakjcBCecbhDSaqqowQvO
UfcCcGhT9YLnh2s7Yc9ar1PKGOLWn5h2HwgcKkbSO/agLWE1SEAwERblGXL4vG6b
0TXy2WbZOl9hrk9BfGo1HxBq7qU9DyPJtHF8/AtKwPfuMYmKKtrssxs7YRoFF0HP
0FWIo8GxsK6UdpRW7f5jWoHQsfea5cURxfNBAzQIYaAW/k8pxqIEgBjYuG9UmoMN
Ps74TwKeGWKjC/Nge8xB1T5470Bu9ab+0yHQ0VJXpziJc98dATdvvOl+xWZfSr9b
a4WjtZqZPoMiiTx4UuObp5M6GrfMmrgvb+ePnlEVkaAajOo0a/xnI2u+euZ5716V
K3pUsBZ3Ik9gaWPlAQ2DBK87MeKCLIswQH0r4PTNCves1c065VQsupckA7AKdUwK
agmlfQ+69SB5+IyrRmWZ0k5VYaGztyzX4Phu4phme7xKw84Q9CjVcUOeu2v5eHlX
lxTx+TPM45iBkStX7+JNQNC/p9djLnDMZc+tRonJsmvNX2+wL9UyorkaqL8O0Yj1
RRQnCSmmANZBKKi1+8HSTw3OJ30NXXObHcEEI1sWCVaabJhMvhfP1yygDE8RLixL
NTxO+mVuDxYCoYs7QyfReg7FBuptjbfuYa4jpcYaA+rSQ0N36RTD4XIZMdldjIjv
aNUzoxXfKrTWMWIIko+JgkS92TFafXvFK95ct4MZwaVr59AtZgoB+ITbeMTl7EMB
+j9duPVX30WnQOR2yxd0eLuAzdScMG4gITWmSEzIJA/j9mYwyXt9gXG4x1BEQYvP
F8lOOLrIFF7mJ54kNQqvBSuDcMLVljj0nllAMBIhEfg08gIhaADx3sywbaAVahgv
3l42FYK+iqSZfLxktn3w5N+w2SOM7i5175luSk8x6XSsd19qcdkYzJnek4448zNB
ZjY+dTxgTb0kJDNMUZGWgawynuubSaGxWxlTlVmqvGvfU6IVDDOYM7o/sWgFYibx
TeEuwEyvO23AbvWYnAAwhzYAIGlPRfOuMbqIPcHICxyYT3Br2pY7GIyoC4fUeQUy
plcRNm3+UgGKsNueIjE75hGJSIz1JstrzACdWa8CJJD17JJvtXNOPUJ64ou094NU
yMNqDCN1jL7a1CVqTCAMJukSAT+Q/wiJL6XE3QbAapkSZKZK9wrDDD9DAmWArmIj
8OrwueiYtdv8Ukq8JieaD70ERdm2vzBJh7Enup+tjKaPObK2/V+DYUWqLKnzxEaf
KZm/QvYyUAQJOx/S0VVg2YDDZBtDQktc79GWrVSzpntTWJxu7Eu1MSMZjlPhXeI1
ENxLCsHqCFLM57IyltJTjaRnAa28H30UWcRn7qLEHZZRFUMgkVpH4bzESMHYaBrZ
jbSmpwAU7mHqh257gpOth5eoi+op2QwVBZfr6qdQvy1uSXnQqN1gvFyVCDaIZ/rP
fhAzzlMFctY+zG6oaWPuDAzpjlkNYvthaMFPJTjHVT4VunIcXzI6PMRx82ZxnAYM
oTPwEhkWtWcXHPejlBx7+99QGnOJ2JyfQp0/6i87Z+/6sXULyhLJ9HkyL03rUcfB
wcsoOBW2ktWW6PUnK/Hwu4krRRs2GC1FAe4rvt8Z0b2EMexy022UzAzQAFzbaHLk
cWxpYBoTouGUH3STBwwUyPEURmid6A8eL8pIlCH/X3cXzZJE6o83S3S8J4egFhzA
rd2bbeQYbx7QswRdAzBUhce+vjqspS3Cqi+iV7ZmSSivgqQe5EMgFkienrQLaPBM
rPXO+FIbNG1QYt9gHklYJnTbK2od2efvFwNsSwk9Lkf7DkGRK7A44k8cllsX1XR2
wNfGu2Tk/OTTpCOJWB8jjm8Mwk0QMv3cx1b+K597/S7AHmoNZWulieLlzUjqdruu
nSSOmwz4zcPGIj+Ag13eXaAEffuFYE52/R89muhLbLMg6CHyy3tEMRrzTJUa9Mmq
q8u3sXsrHkrsZpuMHMC5C/BOaA8As6RypXQcc1xE1zplQkZHT/kTKW5mwD82ZCVn
n2dtFZKFYq9WxSzjI2uSiR4QyOD7uykZI9hp2Dh+p/14HxWgen2rWQKyq+RLgFbq
OJscw0vDoo2/s38t0zZ4yLQ9QiBUg+5xM6VU6n7Ko9JD78zjiYHOqU+9xKzikVul
jj8MOVYNAWXltiEYfbYujPbLUkqphw70w5MtVYQD/AJTjoZwCcsdedUB72ZjZAgn
UhlQerH28/zgFyQw+QN/nlJ2t1z7a6kAJEq2GzO2ptCAHdSOW9tHYpayw8D1NkH5
6KFvFXNq/nuD9K6ZmhbYEHStF8Ly1i4e1UANdqorzxQS2jsiCCPGY0qowBuVcOvq
3m8Rn7aI9hwt2c8Crg2WZWz5yIezKoFLJ7gE6D2uTgXazRUeafmpCl+bL4vmyI7u
EID2D1gm5+QUKiAR04xu3zpMgO5k/fQNmeeBhsNJOtyUDysyy/PGUWfkx47KS4OS
x3nz8rTTzfWZN6Rf5Nv9/RN0Q0E3Cy/YUjB6aO8i5JGSZtfe7BmfqaxjMncuCave
bzKjlMOP+NZC9Hb7KTDk01+B/12T7CFQfCTLj2QLLifWVM+GIFoXSriw3ncFh8ap
xklyAFjOq01lQ24nk2LSTSSqyUFQxfwBmHQi6xXuLvhMsYlXEfS8gNFubeJEuJ67
70EX6wGL10lhxPbk6dlna2GD0BRfPymEtXiOcFQXUbnYK9hgrfsQqzmkND3WoUvL
iiQZCR8MIUfHkLFMS14ud2uzH7oKuYGZA+5VtzrvREcHUjmg8SylcbPG29uIjuHw
MjOXblCsqHdeStDGAGl8yMFAFkMc01/ZSPmAAXxbDbrSmf7G0YGVqj6es0ps14Z6
bDblUziHohYwFAhtUeZ6Zg5JZMkhNQfqkl0XtG3oGzJy4GljoVHhWMblbq4P8Jgh
WXH7NzPorQcvIOueo6FygdGLGVPfkhT/XmUA17n7c1TGZVD5E/XjqTX7vO5v87sQ
vq7Onl4LknO35vnkKHeJONawdk2/pA5Q8Zi1lp52pd614A/OmIL+1vMiIfigUSOd
i9GLkOfCFK6XSKcuVeg4YL+LzH3qPGMxJi4ONe1AXao6TdxvQ/jbP8k5TdYWjmfd
QHlk37D90JpMfaYoVxvS47gVZyBTWsbwOJtENHvEaZHpsdLDXCwmV6ZEKHMi1s+/
rh9Skeyna0yVC4jUg5PxOkkI51m8IcVjxEV9v6Nxq2egcSOJwVhnIAdLqcM4eXOw
XacoFGBUjk6nAIZIYA9FTbUvwlPYhdx2OfeQLnehei/jJ5hbdY55l22uKKWMheBi
3Ab3bvqfCygqiakFJldg8f1gw9ToR5N5uLv435blR10jtmaMINJ/VWiJpacCBUBM
mevTgQGng8D5ju9mfGybdi/qHKDffaLSE49VstKp3uVuVLtj/0vLZgynnGrWDKg4
kFAFtQd4RfVMdpbt/VVPzHAvbyF8s9IT9oAzbPFHoV7jbA1XaZY6fvpb9gnjNVeA
XnksMXlA1E3/xLE+T+ErTqv1BhhbtYWEHWAl35DjMzXwBFtt9SeZ1mE0gp1I00rC
eBvoUkB4ZQDzXgq0QWo6F04BW7PonOjtuWJasksFmlkiKjZJIGZT5Gs50SyzT8WM
2Q6ULQH3M7p4qPO0kHz0H6e7VkHFgIOOD4fMZEsE63JNP/OJpskz+9lx0Gs0rOPd
IC9qz8AMgIdUcWt5Au6wvwGQRwC+q0qIO0R2t7ipqemoBXsAIKVNqobLgS3u2hRD
hEC1jvHuUS60mXUtRZUp4jwWI7x7CjVl29qzZ+eFD+VCHogMnkIeqlgseN7/AfpU
q2RzEQnNIuUSFZSOZg+cJGdPRXUnKbUVhhxKyLfT2EwQsSyTkh7AF57WHTMTglPA
9t0ziu247vn6+rSMD7mhiFQbQNOuYNNiNHDH34LUVZa+ZC0msAIQS33VKzac7eDv
3Zv/h9kSolM2yHl6Y7GxbtzUgodMz2U9uYEwpPNUNOZ4x+M6dLix4rz97jrtokUG
COrjTZtyEr/lRqgXJ8KX8c3bj+Vl/h++/nwzC4Z/n7I4YHOFLtaYqXn/aunRA1MT
ZIzxMFPmsErEtWN0XCtXF1rIVxEoxtQSsTlOvZdiilmDZ95xCF/VCRA4whRjOmzP
Rb8DXlXcXJMuhGtauhgGyW4UJIE61Iy8ZZfYWUOuvDAGxOXC66v0n3YWakdmhc9h
v3OJqxnsL6z5lcMXM6OegWbNcvgs6gotLzjQj7YGP0ZLvxelP+w3R8mH8Bh2GGjt
qeflo2mGQNKJGksyMSRVDkXoyI0U979RrZ1KxfMWfptk+T7lQgl8wRS6q2S5e8XZ
7YYjZu5mqi0KE0QNT3WrmxQ617HdO6Vkohp8L/+FNqEZoeYTv3GNF5W6Rg0kWaj+
ZLL82+w0i/fC15mubEuFRATmlIVjS8cO0YzkFElHo7bV/B2F223LayygvHf5/ZCn
uER1VuU8k3qk5OrxoGHqTqTp4JL1wWKkJUM5Pa3gqFdnq1Ht/fyznphDrK86SvYZ
IEJXoNUnT5P5frI0//v2mbT1lbF3SojsuBjRWn4iobiVZ5gjnsGuUMDzpsXrCMsj
xSOC7743KuvXIXMm+o/WWqHcZGXR44cXq+64otB4B6i5R++/qELmuGUgA424lbqp
uD6nt6ae6GmVo8vXLccRMCtTkRJLvNpZfjaL1dZIiMRB3SgoFPjgtz/SQLs3PhkN
NhyWJB2lbDxNpDIIFKYfP96eO0ZzG0YCj8M8AD8tMUdYzZ6yQP4j9OcUaero1/oT
jqB5OK8NbduOjL9sq4bdu+roKV1frvX38qT/b+HW+3bt0ObAJFaMhuisD7z7WeTh
QBPA2+uPiYFMQjXQef5WivpXCAd81CrVaa949olba8ONQo7jpLW3KL5amjvmboXn
0G8JE/hMTqqyjFGQrp/G8/65B1WnFN+LA8HOKEUOUleDnDB2kuNKBCk0vcVRDyjg
L1J7zc44f+SNfeGM57qTozodzrJazDmzybPilOK1vaGiwUG47SNOv+ya94S62Bdo
oaJDBeSTtf9NX03ohBSIoYgC3fxvHYr8rxgRgYoq2xqQQM1pBn9GFNdc/j3WQIUv
2pNxZ883V+SpH4bneU3SbgMNnyzs41RhLx0u92coDw00VPFccsHu+Ze5r7YBFJUl
yp4qjRq/x5sxrmiXBmxt4966dd59YOWGu5R18CkC91ynNux6CV5fcsujqvjni+bN
rMzjyZOmjVqtXfWdnuwoxF51NuvjBqm+5WqIaghHP9HB0RfKgZLzdSGkFej0ez+J
L+xAFWJEe3kLfZtqLn7q/GYumKB7LLkS8OoeHDNZfhosLe/aF8ppoWVxO6fiWgha
PZLQmkPWxg8MU7QOlfUNI4noOd5fN7W5pBtXIQ1IOPqOxBJuBzgCrqEU5O8U5tB0
os7VYHBx75InFAbOYjAUBBLXwTMkmq2bO6Uag5utgHRm+pTEsssG+y+3EFWyFALz
s0ItEHiNnq82C8dWB4Sh9DX3aDHE+fCrVfmEHU+MqhLMc7/IJeaLM+FQf5iP/OgJ
OIo6WrYJHUr1t5ZWPdniKKv6KrZUe1yTWgMryI4+QaKuMpBz21RX4OtjVEmkoz/C
VD086e19cfvcHqrdSL8lsF2ylHb+CUj3NhITyBE9lzw4VKivin/CE7+wY+XZdDIa
3QhWYC9bkHCgBbZSp2R7P13Zcz6RVD+Q9x/rgePkyIZ/TqseW0g3wsTI+eGyOUdm
NVTEMvdM/XJBV4ilkLupusMoVW65tncMS/X+KNEig+OuutVnSZM3Jg/myKErj8xK
Mtht4LzBCx+noct7ImlIjkwopbqA4VhAtyEzM8BDlsjNJIbDxZDV4Kvkcna7mKxr
x90Qmgdh875TqI5so4//DhfxICT/742ZO/ncsUKS31FN3zW/8cIrgzIhwjRaztyL
edzCD++EnwaTpi3fmJdLH3Ghd3F1WiTp8fBLw4/1e00vtpTsKK1ohFTtXkAHMXk7
VzvgQBzHqM5G0wa0zfdpB5F9sZWgfXxSNR5PhystYjjMqrzWhZ7FNsSeaHCDfjsa
ZPpzreeXpxM3VFWQRLrvlI9e+nNurZcP5/iXKSVD68MV5kWheGx0WCh97xvxgKwe
kuz9M6SSQC4eOm1WW6hdzOuwxf23OB11y6DFYHZ5K5zir0hOP2ffgbVpcn6brjtZ
a3YftmyZ3V7BNbIDR7KfuCJfwJ/Ba1YymvguTSoaVxKoKtSt3MBQI9BSbirfSWD7
euIdqLJWSOq+tyYI9oIXTEaX22Z0agtp9RT/i/JHDuJ0YyjmoH2SJ4sU/pM9uvxn
vpc2LtUBI8Q9yXqwSqyT2TfsEreOBSwkHBnLeR1ioHZSTfiM9wiM4h7EboxKWErH
r3yLQEvTN89qhvnrjaXldX7zg2mxQW1U7kj2P8XPIPCOYN1OXprd35er5hcLiSCJ
fAsgaa3KVWysm0EDfRBFalpDP6ZhEjaQlHYwtlIBSO4pW7a9Qxqf2XxUUrO+NYLX
iDE1niEN/V7eT6vGjF8Ay5KYBH/03lmaO60zBQ+ppjZR6kkoiBbs7c1ggGndHv05
wbKCRnmu3/JN3FVuPfdBLTqoEKjGeTtKGGr5XgRqmJVpxsIfy4ptCLL8iS8ZRMIv
Hih+DJCd1WrXSTIhJGCpRY0Is+2mJoy2LK1opjDMQhs2LuPBv0A6Maq4Xcf5xGYe
qOTK+/exKsfmclvYYxMoDv5D2q05GvATmNO2Ht4a3Pdb+sZ8qsV7gDpdY3uSastA
JEMx/GpYRNklIuGjPu+FFaCx9XoiQ2Fytj9eb4/jefaksN4x5R663+vVN+56K0ui
lGl5Koj5SuIQ8dmI9Hqse106J8c/xej2XmWYFLx6g7cjOdtc5MG+rICE1muhqzwr
/1f5a8mUi1hIc+/Vn0sonuWKGq7+AQ+OgC0U5I+xoQCjYFo+RgvQxyjf2yYL9wug
vvqkB12L+QzljLJ/Xzn0aacVQ1u8UVyG2CFhsExQaebBCQTHsisAA28+xwyOS3eK
BT8ERHQI7xQMekQBBATP+DXt0ZvAi7EpghpYKhuXeJEdM6tHSKvWEydNf+Ye9jIP
CVCrfZ6XXOlDa9AOLVJRVeRaWEej+9jsLgHjZAqfl+FzGh5q6D1Q5j0UmrZ7Y7fB
ilaXb1j5ZzTsUAOCMSooV7hTza0mgG/g3iVOHyCpfxUeJ04hI2dFpr3WiEG4TEOb
TYqP6Jp8XMU7I9na76AZQiHxLUsJCFxaPtsHpuVFtIPPfmg8IO7R5uPYBpLwNd+L
yn8Q3xCmeDQYMjzN4qA7ist+R4jcqhI62Z9+CPdm+hjWIEMtkNUjIo1Cr6AqIiES
OVoUdhUwMHdAkeNw+0+oDAsgk1nUwZS/Oi7kWKosqxt+PdAHd7EL52G/jYdEXUX8
3RiUPNV5uurPwNtBEqxm4tAs13v4eNfv9DS7r2u+MBQTjUgjNMDRAYbZEhZSusP8
4bYNoMvEt12056800vN9dgSdFFkRSIEc+SKo+8uaeB5xm+hnTqz6IYxDcA8WD0Kb
NYTJs2ip776opU7VZdBJsCWtqaKROCTaYHMA8HKQvkcpZrALfcq0mQWWw7XuFtAm
l5mPMGe0LPMAKq6JLo6diUYAe6v3YBJmHUiFnI95HyrAYFXnYEjVOg6iLktZ4ujV
ynnHC5SnowQ2VAWoLsNO/CC4TPnSh7NbxpCrhoklIq+LzcAa/mvaBv03/xsTP+6o
an6a/lGKeabtlexkyOOhcxmwlZyULlEErfdj2yxhcswpqN1PRa+9o++e8Xm4gF7o
eJWedgHyFpp3bbPjTjvu7ABlOlT1JBV1zDh3+HjGXDXGPgtm0ndtKrx6/FvhqYHL
WYILv4AcZFHUtpDXbfzU2iZoVAzK3RsGiQqfkEnUOLpnF3kpspKdTchbdv8GzOkK
BxrXN7JY86MCfoI/F3P8Ng+ImYD2GJ7ygBJMxTV+bBRUk/m1E3sQKkqqBi+8vvw0
rsvq0UdO3KVcI/w8HuXzHzSNqXhNBzVlIex5PP9WJYRP7YcStJuh0Iys2aIblHV9
uPIeAYUZzuZUpDXnIsoucwp9yJ3oY/O6Wm1yCAKpx8nIWNEbJ3O7JGTLJpnQkdUL
PlQosJl7VpXQKifsMJkT/5dRGwkV2FwoOAwspfdMvs6Xv18lxTRGBXxOgABGn0rH
+VkJUvALaf44Cqgka9wqxQX2990wVbmOJH6JBTqV3fIQ45zjUM0OlvfiKR0ZLaPg
nFr9mZ0XEx0sZ6CCupuYs3sTf/qvcvkKfPkq2gw7xK8CKjdq/Z1SCAkj7VKKGy6l
C9GKZL0FEXQ8Ksv1CAIqL27UV407CGNbVwIr4PEls8OGx+BdZth3HMbNk3rA013m
J5PKgPi9Dg+vndm2iqFPZteewXAlg28XG0bCXQcNnpde1f35o8G0+WZujfi3aOSy
9+6XvF09ScVCKw/bnCpdUMcKoDPBaabHlMiCU3iAKvYW17wOQB7hcF2VbnG8gTZR
nplq2ATA9LYplwlrWFiVRydl9HZcK3NXLeTfn76C0czor7w0zoQBmZWpyRrmtYGO
6Y97Nppl9lL9+H4IsXYURfkczzFHyEuhQr3SWDglhPA9QzPcLN0R5rI+8jd5riuv
4nk1/wXD/4weH5zzwREJzhnqLzjHQ6/MIze3ZZW9eM874HHxqalhzhPYxzlMisDm
Z9TI7duu3xPPv3y/fS2RNtCqOLWBrk/85heDEjRC8umNphJ/GqdqqyuDxAFMzeX/
F14rTT7lQpWKK/dPiUSMMjBGWaHUAFAoHX/by3ZjzNarZsiYYZAxUHWtKO7Jxob8
suJkVLEBxxGpsjnt4XV2ltfnlsHWFcWUb99XsVnYBaq6odcHB+dNUHuwnlH3p1bS
3VUw9Vxu/kDQA4qGuYW4lo8D34zbDGz5BQF+eM6Y5497qLFrVZCe6vpT6xL5ES+Z
NnOLJBgBwHG5e4Im11eNFvCmUXIjIRhFR5nMpCrFzeTtLZRL+kiTmrkEuKued5SZ
PQCMrGs1uOKC6EJGJsTddPKbOIzroK6s2r6otFN3uQcs8RLOHXGB3GdKskWglL79
a1mwB2HZVbfxvYmwax6NnO2FLpN4rMGGTTHLXtFrJK814MmOe72KJuPmcTExYGbT
5UVAEvVmn1OCQRI09AH8voKiP0HemoSOjQlmeVtazPKweC7y5+w+bnmA87kND51k
kAsU2EqcI5uEdBcvVtf0n+UrjdZGn+ulVt2p2FvdFq6X58KDpd0+h7YgXD2CrvZh
cLRrms1/9H1M/KfQeRwjh7zp2BgTF7PpzhG8T9cwLP2mSMK/4qnmTceQvY3yNToK
bwW8n+HYyYhSIFbnfBvY+rXsjHqnXnLqbstg0QJEa/C24soXeQVboGcU75kLvv7b
7T4LBt15R/OcBHggflji+ea6YNpQV2r6vywfk+TSxQzg68KA8CStJG/qDm3yr3oX
92ufvuPpQlxf3+OkDYXdXqyVP1lbwCMTju9yP3kLalspeNO7B4eymZwx7CQ6AEmS
dsBM8bAW1gvIb1KFSZmIcsW1nmMiouNBLV9HzeLN8CaAeurIJdwqCpiPAmBbBh99
xXoWIqi5Eyt7qRp1RfWD9Nx3sibDOXLrlXmb65uZKP1QB8lYKCGKoTdslwmFCcrp
2PHbEy8KmfcLv3o0i5A2b0+Vwg2J1wkB3voHKNMxa1NfBzgU5QKOwmP2TnBkqNIe
QgstUn4H3cTTa2bZ5BSLytG6EEkNmRXkAvOxx/kChoYedLvpcyeujnPm2Kh1IJfV
e7mC9ZFa/1BEl1hoojfQc0GfJ2VvA3NtqXCHlUf4NpK1vIl4MCcxz0UfDMhszqma
lh13MgWpd7wfSdoa+bj3IXL1g9eVmbcUuT9Z6mtLkhOMM6aPyk3WFl0OL0dDxot1
Qnhw3BkbDtJPHDlJPhsqQ2ealK/XF2fY/lWJ0uhcZE/bY8eRJCNqudI5onqZUlCj
LTiD16SqSjsaTc+Y5JxI9pqeME+gNxKFAOaop3m1tNfd8COrfHfQrhxnKPcPLHzx
gOcQhUmRQj+kamAWad1IcrDsoQUFbgENUFHvLBHarVBzqsqU7k0OS0fE7sjzbmOV
2+kDBSVnQk2mrLd/9tIoJwLb/Qp7fXaMwdiO5if7YsKmeKW8IdpJETLlI7Nc/oeb
SD83qc1MhWp1LATRKtPASCRwNCoYAz+NPLLvKF4qLMSqlNgBr1yZ/P5tVsFspkng
S8dIn3DwJiNT6Nsbc5mEqTWVZzrKQlGerSNqas818qqYCG7U9/3Wk0PfnmO5wVKE
N5a2kiumoFHzzxyOn5jgrToY8VkO2JwP1AltOhWFqA17VTtPuxmCsDkVfr4R70fK
7spa1wHAFEGj/jFdVRTxg9sxcgdwGGo6at89TKt+JONvx7/in2IMNKyyczqSR9+F
/4lPllOerAe6JkMQLHkpDv7pRmSSPf3wWexrxHYIlCs0G3OMShOeTZnr/t8o+KQX
o8Ad8UjtrTjda9Y0h6qMc4s5ynwfUOZ8DFD4lMOXSyA+8JYQCUs+nbgneI84DnJw
ujLCPKvTWatdWpg3UalV+uwuAlxbiFHOow9zK9o7rL/IMizi1TByEThFQAqMYrer
nkds1qA885RJOHq76ELRkewzcoI0qln/8xJYNbUFS0jxeeDIyGAlLOlp2GCgX8YN
XsF5z4Z0+6nUj+45XvOq2o5zi192E0r7j8/7l0M94t2J526aB01UESa8tV75Tfmy
6Hcrf6Ecj68b10B96O6WzaB91SXqsRHtECvfGr27qWL+o+ZiWUMo4A0ASiAB/wEc
eTs1jflHl87jpYcuuRN13aPJLce8/xLujGxJKVYenvQ0YWrwM2HiZMWsPENjpLHV
/j7CzcKVHUvRjcUFTEeuREiFLkWB+q1ld5UMMoDplHL1rHwdnO5nL0pULq4ET4sv
CATdsDrAqKrLomsFRHoeIByi73nurIFIqG6VbxfZtLjxr1IH1a6tK8YWm3y5mzYs
+N353dPVFbZEWfoJ2kXS8kbpFfK/um+upY1L1POj7d4gKzX30C2oFRygIRStcSm8
XJje+YGPlc55hbHzkIePBbxCPpcE69W38d7EyBTXrjNH/7pwbEgBVDuwiRn6X3eC
iBZg8FPnfraTaC8WrBnsdi8ZPJ29s8T0/KEpUpRKeIzawiVeqTxqnUsTujLTEJxA
0d5afZZCdW2vGdPB+i4I0O4JmGOJkXxwq2tPlyiskz0dao20wzgAjGY9Fxm44q9q
296s165JKtOAB0SiiMyr4KeeiwBbSTDI49DxUOG2vTPryTJFZwTyoOunxE7UIwfA
mdgnyvc8/JXQ7uPVMkRU/CGfKJRxMraI9ZkKnxjJiP3Lqr8Ny2xAABIKXsAal1BI
I4zKOI5KclikUdhwtl5BlhS6MCBhdBCTeCHaIEqhdFjcFBrXkl8U7JUdpnkK5CEW
A3DHj13YJyRFF+/fDV7E4sDNG/dmoewErgBj0pZb46E0t0WX7QfBfzMM6N1jTZ3Q
vEn8PNnMtu9bdE4RphHOL2QdnRaJq5F6I4QofM01r1tRe3lK5bVVszCAzlYN9Oba
mr9zzUmmmxexpnGPAH+q+MX1PsMTmRkT/o6etx65svdJd/+gYCCSbQEpf9EJdMgN
K4Cw36O9ffRXLPA9AOD0i8R7ktDwlFzuTfnNPr17CJbpSJuDd2yI8WTmzhQlvAxB
B8OLvE/hb8YaZ1xA42DG3kUJloMtSn0v0R3r+FUZtGNVUILhvqBcm+N6bvw9Wxlu
408NHhCGDwmjku6Pad1LNCyCdIO3xY9rkO5xI/Ov6LCztyX/t8XoXDKi4fsi2obM
bJ9SBPh47GtLjS911QA1KkHYVShNNcFO4ScjWT6vQrvGi2RYOrJKPWE2QxA9c4gJ
tRp8QLXC7DD6K1bfQB+pz1lyVC32AFGOf+OuQs6F75sa+fuWLp3xWsHQLNZMZSd2
XTOJaLpzeNNZyLF3LEHy8hNsGnw/X3jnyYzK4R7Vv6uoiCQzE+OWEAre6AGOaVOs
yiIYAP2/EJQWdBTwOltPJpFZFaNzHSHl5lfV4HNfPMPtp/Z6hFNUTQFHuQXhPq7G
N8dLjTsagvRTWr9ntuj+qBbSCWvTbTqW+wpyeoyXFJZ/OjyXIfGSXk3/7VWPeEq+
JU8jkdJ//4yMy6xrSu8+lD96O1vBWxdoLub7GzjsxbP0pGS9uHLIVgOInJowO1PM
jY/Ie5/7MGbgS/8B8/ej3iu91pLQgo6E854kMph1qm8dNtIEyOuHceocUYBS4m5c
lp6Y9vV4P2o3jrbs7sdekUyjLYuSKS5T+qi6NeHMVAvXH14+ZBkzpZnHVCAipkoS
yoqJe4UvcEWcNkc8VnetP3d8i7iX7Fhy9W7jeE7HcHC7vMSeEFdi9BCrDyQlOWz2
uyXFkr6WW+eMKm25XQEP3/W7Gb/ALw5YJWc/hAbJcDHO+6HGdcwOKYmxMzrYPZ7x
qGmEFcnBHpdDcEd4YeFXjn9fLJPck1MqoKoHdFLIDwS+KThAsOD5UYZGzTsc9e9T
YAAWlNdXwCQQjhVSSzHEzoQxJaLfdvpvtWBiuTlhUadJGj4esdw8JM1kMPJGH+je
nAiU8MkSZOMij+vLgnZQf7AO2zu1OyxX6EC8tMkMcO8FdQWwsVxRSKr60kgqXlS4
8FVYPAf6OsNI39rj0AHeotD9DeNacDaajRNN+83KWrhre7SmE4+So6nmU/uKiZ+k
tpFEChr5Mg73B1nDWRXbZSgWqIhS5kXD34MIpkfXva4415qRBYKaaMFMc2l//jyZ
kgcG1uqdA9EiKTg53ZXhBzDQJ/QuyTO0vZBJ0TJOZv1nZsJ8DTYpXCwKGyE3QHe4
t5UHTpqTPYBlcLAWUaWdMwLr3+rUWx/3NA7pjwMNdx413NBT9SfNc7s6ihx0n2zr
ZC3SHmoMkdeZF6tpSZBJl5dzqnzPQSZxT8/aAXvY0LrU5drvuF/Usw80a9Q9My1G
IdwbmmTblq20q4c1OYRITpzOLvh2dDu2QgffqdWy4ctdE+JfV9ebh3aMgDIu1o0C
/pdqaod+FnTiTvgd6uLUCWK7SfL9JCOCssoeCwM31Hf7lM5nWNTjeBu3r0GQMapd
zW/Gu3Gq3/L+7h6xUWE7nzWW+srJx+Pb2lW/kaDgfNU5B2hsZxD9MTF/8NL9Wft8
oAbo4lswg4INQCOUZX4KY0SiiP+nL3Und+IBxMhJnoBtzuERGj3aFAMFzZNQ2d6m
iL8w7FpzeQu30bwdtikQW4pwvPEMaHxg9F0sUlknuhbScAZIbiDLKwOSWBNXHLxX
UUELa/54JA+ZOOBQgcR3xKt8H2zribHwrncteO99oeO80eHE0dvibB7G2fJf56H7
GKYzHTr3z0Nn2fOjY4bOr/dSbEygsa0tuJcFIp8BzlLPALscAZXgbmzdzRnUIiis
qAto2tQAAXhiMBEcWmxnv0o1mMuWk8+fhAZAINTUqaGTczpEpLyk5AGQ2BDaFTwa
NjR3g9M8TdwdsCCB4NeZrAsJcyuyEXL94u1Ys1xub1rNKqIjxpGS/K8ySe1DbjjU
cIqYPhhnEXZpcmK7QDdAcyrtSS8LtR2rO6YVi7gWQIUdYRhVhkZ+FWKcN+LIfZVj
czzgYMxADcujJZkVoic/jBRMUcfuKfKB6t5ndkL6wEaw7Cqu8/1Nz0P15VHKzkkw
yOXbmdXe7G1fbdmdjxdVMjZcWjAEMOab/5yAKWU1GMTrGHyiifKLWmZQZlEw9Fzj
S8lAXfUybiDZtz8YXCIEr4XhwmNdQPcPusdi3HhIPBIuYMDZfstY01rp354/XPll
4sESXYi4etAdImC52gg3AIIvFeE9ZYiePauF9fkK4FqHgdUPT0gzw6+7yFVR0IWb
vN2R2tWAcfTDh/NlBxuTUS6LfLEEXwDLiWohwiONXfi9M6JLaVg/CMTQfae/f5e4
lgbBOAlwjaLU2sVlCw2z+2vRmRoc6bSL3VKjYdJkFIjm4LH+QogNs1ZfNPDvd7it
ILLWY+b//CIsQiejybuqU5LAE+omoitflet+zeiEWmPZUpSLAz+wXyoDGqJ1N8cR
A8R8wVksQ8sYZkBeuVdMuhlIQXiJPQYKlo28HlBezR5FtFfPzCBMd1rfK747cHrf
2pI0zQOCTcY+ZnMy68dQThgv5LLlMUIuVDjXwWf90mf/+KOa7AUsMnkcpau8ZLk4
X/ViKTjgN3Nfsc+9eoVMXoStEszlTniSfrOUZlucaFcrCQkJ6vXwtP6EbcCHxUs0
8IiFatrKXCc8iJgmiI4x4rXBejBigiDV+pPM9TpsMy58zsAEC1F5qPDMIfgkrUCL
7sLkEzmuajmWxZR/YIVi1gstH6inVs7AZ/XXiCfWi4Y1LqM/6be4YLiHPFKFSvuS
Qc/5w32ICJyu5PD8fNvr9jpy9wUhzdt2e2pFgyt6hsvD4n3aUHZmm259r/o0Hzjl
+i1xSMNjPMTAEJTEN9qBrXhq6rO9yoZvp3xpmBvAFkVBpjRqsrdLhOYWAb5QtrMW
/9OoJbS+upnUDr3eiVBLeThbQS1wx+FiquE7fNnRcy0pOXUWUjqYljSOztnVylIU
PbX598R3H3y1YB39jq9bi1+mwh3xT3XOuzScP6QkjyCAltoFa/ygVB81TMTVST6A
hGmqG01twLn6l1w0zXPmHePKCX5UjPIgdcRYa4gJjIKP9ov1BSs2k+EgqD27LAcy
xwSuCIr5D6HNISbqowHtCZGPHF/1UnGRpYtrBG2AynMWgmH10UOv07gShVKdjqRa
Zgrle4W50UjmJGsSNsBXusBpJ7KpQUPxnModuXPc1+V3Xe0QqyUsX+gyX4F0geOx
RbskN7XR68eSBx7LFpV9/AvnJ2ZnN4TU3FxsrqZcEkvA7bKxEAkdRcKNTgt31+29
NGvgIiR6/xkEHrXVIsDYd9fxEhKIwybKlByyPH75g5sIuqeJsV2Fo5VsQXWRw53o
r1VgfAcXT+Ex4JVZKzkk53yfsWUb4jIWxgz+HVMHe+3QgQ9NtL2AEq3Wva0Ni94u
BTqgs8GQxkTAuxXCX+PDk+M+ZRmsSqbZORCDAzFJFrEYknPXCrb5FGpa0CfTI8qI
rNQ7iAhqgdYRvhFylFqIiTWn6vzJ9hAaiOre2JtkYFL1cnZ84nh1UL+Esm0TALfD
1R4IyQySu9L3J8vKvH31QnfgoARSOmi4gaNPTf9a7o26UoiLvx6aQ6HrN+tgGU0o
/mjg++YOlCtZCkUCZSL8VAAM7tgEs2MhG0j5WYSoTRLpM0M3+28ma+AtWcb5rGO2
9AhkI2PFDtm/71M13hS4P70aWvUR3DS8QICbJlyVXG1qxr8c/P7awCBUk5BPEmZx
1I4k386ZXljogQDFSUl+ColvaV2bS3DAsaGdrGZSHk2OPRO2Pp0o1dWNRO0foKKY
p4SMmx3Fg5Wcvrf02CAJWzvOoRHOLbVTToUeFM/jnEEP2SX8Tn7Hj/BS05qlG9s6
dlSl/WEJLJKj7CpAhaqgUMTQFamSe7gtgFxgT+RruKe9DR8jlk/8ZIcuNiUahCJ9
vdoMKepnIdzxTy2sae9PYC7O15HHqflnlQ9JvbBSFUL8BzUnsK5W160YYUB2U/9A
5omPOJ31XiRUGnX0eCA0EwKlQNkKgNYvFHnME4n8jysT6nc8hi12/bHPd1UgSsTk
HzFk1yd998pTs+3LlcCvYACLya6uI8rjbE3cuzVIosQKjSN1lfYYx2QqkgKMfBs3
vbAOdbzcV/dXz5LzNeIHdiuS8RxYyrko80AwDP74AeE5x9yoBCtKkgaQuTIZesZW
Ql5X7lWu2uwCEBzVTnkqNN0PGYyy4MD9kQ5oTTRcWotj5IxLyBqI0YtLCq5LXggd
wj+4KezHF548b4Sd/g/m1iXBEbPVbvjoFTA+pxkzgBKupJPvHakE2fpmEgGW6t/a
TO+5HujEn4k2EsR3KvemQT0WD5X49Auli4PuuF4VsvBme84BZyuijMdz1fVdl+6g
J0qYfiiW3+y2VT9bJxWwNfmZCKS+24xFsllKcX4RUicHsXw057VsRGtN4WYCXPOJ
bKPhyyZ6cR3W1pnwvm+8gHrOQJciqeowC5TzXcN2/bdClQqBOZ/uEr3OLHntDDs6
YIkXjJpnQ2XfYpfa5cfJI8aBywrue5FAssVSzbBPhexysWLN1df/BhdEC3bRA00h
yXPfKw+Ir1LE/fqw/sTq2jznjLrHHZrLUlSf/tPoIiiQR8E9MfF8Nvst/+o8kuUH
80phrJ6aXx+eOfUGD487Hj0tJiLGdNUHan0nukBGyouE9vnXSfhxofn3MfYRxrwW
jEGIgd7klp0N+HgyZi34zu3BTd4CcWWKOAH4cfcAtU7YiA8gLrdvXD7uFnb3zejy
DgyrwpgvOWvKAY5NJzV8gvFN9kVRs4jJ7xeQ9uikkML2fDjnz5LUbpCVPVH3bq3J
lo1qIIPV1A+DGJHBwd/VVJyYpiGdhf2IxTdOKw1hCEjUrQ25iCLDG8F+UgyNDXku
uUKPyktYU1kSXkdyecX8fHfVtFmT1dzNaGSr9BItkDbx5UbLvQpa6oCOZF9KPIlO
X919RykZEOOR1W3FBld/QMKsffj/HbvKsxllvuh7jlcg86seSPgh2/WqgPg9XF0X
MfymTBZ5QA4YmqIpNHQUzJVkVqzcQXLrLCS8+mEUts0Ycxm5xiKrpQUY3y7FfHTH
E+oz69XqbPpxUqrHHo8Pn7dpGh5jtsp7FcawNpRU7EUoteoji5RUwefx/BBptwgj
1bWcyNABFqxI+rFhzQhyIsGDbEjJLxuDZ0WpnRIENGPQpigW3E6sQTm8bcmJ1pWD
3HneCx98dY/UvpbH8ib+Tihl4Bper9o86oukG3X5ZlP0MtOzqJG9NUxmZpSQuInf
p4wqFBHRAI2kgnlcEvm3Nu0D+KWpDp6o6DRWna6b0Hja3d/Iv1jGCsK7TvskJI9z
0iaGi+Z7dZe/6mS/GEzQF4a/iJBSD4gOxXQOjeCLi8Q4IdoQdE9YYralrhNTSLHT
P2W0j5hU4jujuwsDXS2DjWHtSezL9Z21XBy8f60Z5fCiCAvc2rM6tn++LnevboXF
P+fAAgcO8KW5tfYp5rHjjuUSLmOGHCCa2Gi+/C9Zgd86X/mWAUGYB0kFsW9Qg1Io
VZs67NRncERP+Df5pC/lEA2zYhRWXUZKmqiR7Py6JnEW/756CaGZaIysYiIE+UcE
iajJ85jAEkx9hBNFBINgjdXy6BAFqnPR3X+T5CTan6PImbZ+qJbhEd5vhqukNHGG
ANWyBm82FG8cM1A6AN6IUYN+ccOewUgabmDr+nofA/0G4WXzedL7ywKkP/smhJLX
vvBws2fexs3HLDszHanBF6WrLfyNmMqYUye2+ostFzlHQWvCiHBTnZHdg5XubfL5
R0hxvLZKo8ERMCXmDWCLDVo6fgGyXlsuKDOwPxQ55KPkOKoSrdn9RZTBug6dM51y
S/aW3Kx4htZJtxPl+ntXCMgmR7mr09d7iwtturv1L3S6igLbfEQGp0/YKoYxxuQZ
7aNp+ecGHKroQTmOIYNd0122o7vIckr41Pto7sNElUBNrJrVa0Nje3jZIuBqXjO3
5t2BJ73KCKHKJn6S3FtB+RGfoik+lFmDXtWQvkGp1ao0uwx7AD+0nyzYjkZkJMsk
C5f28zJN6RYTQeuvKvGlJKhCZItMQtIiXlRTU07CFAoYINpgEYMc+QROg4hIDvmf
dcI4Cqjxb3vZbziIHkXcSPYeZFb0LiXwGy7hRlr55KF0m+UuDnDqJRdIHLa/U73c
qQvcC6ofyssje0iqwxLFt646MSi5K7wZp1zxyn01Aheb274IMSau4BL0xylUuN1l
x7UX2BgJwvUeg8h6E/vzkHrrT7X4A15t3DjrGXG1oQVzBdcyDzUe1Ylv3QLZ+0Hy
cuCLk12uZnyDJS1JyZjBF4/wHRSt2Js+Ew+RUvpt/z2g07EOoXHrdh+YR94EQ4Aq
NoLnYgxfjKR2KixAUeTqgZFW53akXz/N/4opsYlNGtiGychGMOxeCiBjWWKk/xJY
er6KbsFKy+HSVzcYENVKuptbd/mNs3VCD3TWT8U9ttMB6Hty4nBuGRyh/Nxf+agd
gt6PXRdhOJOmDbncCXe/0WaGRfeNJr7MZeW0F4Sf+kHvsGgaq3yvgNLYB88EDAfD
s1qrtlA/Zd4R1zAR7jMUVx7RE9zrXAjlV0dUD6iJ52TCbnSThosqc0F1Vo74LZg8
6tqfxQwmV6k9QyBnbXN4BG8MfiZ2BzJ6wUgdt1su1Dw5T0CkGCjWQ06NI5Obs5bM
nSjE3Rc0kDImayeRjJ9CVbQKuPw+MhQOW9n8ZSaV96jU5CAl+0xxtjcFAva9jhFJ
pIu5gKydfV/zWmL/xsrcEvvlxgJzIVFqxjfcx5w0Qqyj/aTbaQrdogsZHWhh2NnC
vgM4aVC8hucERAgOibE/Rhdiv+y15HXLFhmu2zM+KJVBvNTOZKvGv8SpN0HFOInS
f4snTny2kyEFoonDeL3hCCb2j7NzoMfKDoLnIiBAj3iT0jP1s/tQ7O82HXwFG0NI
HbVBM9fWvXZWdQsWN+e8nrnz0t277DTc4JcSKt4HGj1oT4afwXlnbyPXHKuLQTSr
kfW8wNcCIbeEyNWKtQWqFF/QzZw7fDFMr2/CKr0d/kiy4dzVlHouGupYAp4s8ukp
oYIQGqChK2eDFR6WY2AMDglTKq4YC8DwNhzfHDfkoN4zil4140v2boGCMCQFm3KN
9IMdvg6cdYoDtfD9Tq19ve967p5vjqJfvrj6RbUuK5c4rOqe0Se3gB+K8whHDcSZ
hd7TNiI3cTdJukphuSfTuHxhqQDT3KJBDQ6ZiPUwb7Wn9wG/UKnLlTOpZX/IjxsO
EB29UhPLWUp40utrQ+xhnTlaNt2aixHpiW4n4P1QbQiqXSLx4NlYX3eTDtu5yVHv
NKdO4KtSL20FS9aRgXoZW8twti4FCHDb9HzHsdkirJJfgpWWP1BWE72FA6pp2gAc
/vwGsgh1UmRFWnzLXYj7u+0oxddexaDF8Q2AZ27eyRjngcJwoD0zgzjkb703f9GR
v7Lx8FaLfYJ6OXQFqHCNY9ovFSm8Z31oLJX1Q0V9lPl2AHtwDNWlSnzWfuDFQUXL
UJoP1vYUVpLlNn4eNavegmQkCjsz8bOU21mpU1TIeBIuEwFpHHceTIgky5mojRcH
FG04oGyjgQKQv1J3n6dGf1U6AbnyaCkgKr1vV0e4dxp6vYGx+gV0osB70wav9Awb
Q1F1VyKKPJkihWFetTCR7nfE4tkjdRo5HxuTl9aIqqJ4M/EzqYFmWqn8NBmxIl73
jNhqWrwkI7y4MeNapvQIE8I0HDDJfaX7C0+5M+8+yfNyxP/H2ltUWpgnPEeTxStd
dhnR5odinl2pTuguXgcz7Iauhu9/m+7Y5vm300Znd47sxv+u86G1ND0cYvHcVbbi
cujeLjGNM/0HAI8h5bGUIB0tcdrzhmQJKvVJkdRxIq0KYpVRSSoc9ngVQZN0DnZm
OavjfgMbpM0Mu2agmbh573ZkqsuxfUqK14eycvxc5umL/bc8PPwD+WCt+ebgeVyt
1sPxqSNqQOSArC64lSOkM7AT4u/VezUFC6bPoGGPaKmza8Z94dPG3Xp48l0+XPJV
0SgXk+YCW72vCVari0DGnC6YivdF1mVWVaPaKfsDO7uFvsQu5bQiZyJvSPj1e3wV
stzCHJ1ITayJg3tBzuPVmmU89h2tAl539sF65Dy9E1twKFyWh3jYys44UyXNGbLz
y1W2W578//pvoe4/GbOUvJHCgDpEwvze+IGI64+D0rsOVQrTVrT3VBTKQqp2e+Io
nzWurXqYn0c7Ty76u6P0Wr+9UEHhXNFHzUDIsYUMkSkBUYdYHQql9joUB3QdAbHQ
3EPbjQ2/+DkWPe2a3sef3dEt0uuDSg/RQvwWGnnBG7JEsadvgxSFf0apxKha+I+3
s1F3deYOumqyFUiYWIpvzfERagrBzi58PlxcemV8Zzo5zhE2WsT1OH3bWBaFEXRy
6p70lDIA4kcIYLjRzJ6MmjN0FNy0y7jR8v2Ox1St+jGWtvKyiVzm8U44SnDShTGi
CEYQC+xQ7SEwpUosQ25bZLqpKoGyGJ0lMpw0i9Wt1tIpg+pkNu233MDPgfE8a263
4WKFmMw02ibP5wOWULqDTLkeZBuCs0wih1pWY+gpOK2i/qso3762YvhIH95OtT6k
Rnrg3ehTgNAO1gWSc4w0Nuwc8qACpfPrnriqNZ8K64JAFmKaUiWzfYolTugpHbs5
bQneqkn8qm7HVAeMMIggBuSsQqX5VbU7taM0Rc5SXvGflfNKhp+YKISlRaVz2fLq
72F8V1rScaZGvCeucUKAYlnTmKxKaz16kudkOJP8Q6tmuMU0JCesW8Mf+ZfEd1uo
x+WpVYq+Msu0PSZWSDq5tw4ZDfVgMdlNUqGK53w0y2xJMOnuh7TZimjP/kDLzQbQ
cgBAR5u6AiepB6stS6hnnDfvMqnFptiE3q/JL7YVZGeX+R2BVwpP6k8yA4RdBNmz
yj1/+Jbk/i/CH1gjh1QrIxEuMfK2CiHoC4ciHlHqWpJDg8rAw3Vkely8+Erii3yQ
+7iBU/PDFvOCpesKqTOpej5wzj5FWqNlNGS3Bke74ID/FNe0eV88u519moIkGTZP
JwxXvrUUO5HR3UD6Xl5PsBq2D/vmHQkD3FKllr4Mu1XgVPdGlswenrPL/66IcXPq
FsEgv4Lvem6sEaxiCwm9iDtPGqv2yoU45EE0IV6qtmeZTKgK+cUaNJLeiJd9pWys
Cw1f4HJgzACyK/DxcoKqqEpRj+wJwnHc2ftBHZGRNUUylXTJYQ47gVLvOQac9VTx
SPrgBvEmOmNw+6gDZHPLtrn/+ab6fh2kwI6Sf+/2qlYvZf+zwQaNDVYszJhqiLff
KyOD2Lbaz5b/AMOmcKelJIB1K5zPdmu+uvkOTk6GJfLsJE0d1g+63XHDlpKoOQM9
EqfzIWnOMR1BPLnQGc22cxgI/xr+bTEEaomrzzy9HKYmoHAviNffgzzrGChDILpY
dvaYqqbyxTen8E61sygxwYBDp3BGoWhu841Ngp3gWbuQGnetu8LbZISJnpCf3ck/
n6IsCIEMapuX0ClBoqcZVt7aXlWIIwCoOPgUUtT811HbRHrW3ggE7GJ+4F9j6Mjp
8ggMTbgb85XvXZd2fHM4hLsTjkFpuz1bJ4ncxgfugYYySyeEr8wyVxU6zjpt2IGq
2qdUFnYg1v9+LHSNg/vk58vx12a6nH8/ict43+bn76oGbmJ7WMTEt3fvLun+V7tk
6iz4WqFQ8e1BBMAddBF3dojWYk4iFGVWUlYbYJyE67sh3YS2mHv6OY5T55TCjhNj
58oj3iA2W3OHQGDE5feevbgc8FuL3Yyu4nnlAfW/HR1UlamB1BXgsFYVAvL0i7XY
crsS6hukOEa48GPyn6tUkjR9eMHrrECj3Y769Sq0xFupSGR8dyLGtzklRGBPL2W6
N0Q98ozcI8B254M1kXd+41TrMvqLodbdRY0kLku5v9MH4K4fAsF+P3N+cxCgTg1U
RJSKaOI6tLOD3kDa6kjCNmIl5mxRdiUT2M9Q1rMcftphqPp/9vnrhRiGd+K5x+vb
lef2kjrV56nH0ZNNevbCv0BEDwzM04c7z1mXmoL96MRroN5im+/qo0DcPhGtGXQN
PLzvrxi3nJFI5Hz8xO/oeH8ur5Tqw/nWLaXt8i2/767teWdvpZ4+zvqXblJlqeWC
o0rRH3AG1d6qf05ExpE0o/YMJPA8xhIMZzbcSVsczLeRsMTTl94WTic5y5z//gB0
DAfyngSeuHYCEG1AN1oVEqVQkpYeaA+dN22bZLIZXN7FDqFdWuNM2h50+uaLR0ZL
6PvwY65cKDauBFdVKaXiK4jvdIn1vbVUvD6Hw56WcugRdrazj5+vRzhBs62auzVf
b+kK0VQnq0ju28MNEy5O65dDll1tYG5h2z/0OVDBzMNgZBWvew0GMwgMsiYcwjh1
JuKJ0kHX7Z6Ryr3/stcGFa1WQhgBEb5nZJdKCE5hk83EwyJSDkTm3+c4JafQ5rpG
2pH2NCBXgbpc+Rc0k/sPpj8q0iC2JJfpDcdr53E73I6MCxvn3hEvLCPM6IG8+jew
u57kcRlgvii1h5BFPBeap67SHNu0tyPrYuUD2ps7+LMrGTSDrjXYTfqV4RTeJYZv
/SW7KDOwemgtZR65XmwJTgQErB+I+OhalD5bBOzbpfQD+gldTm9aJIXfOVLZ4Nji
F7GyNuyjo+taV7fqG/l4pCTtBOtGbjANTkv+ipn6Uwm2e6ZIaXnf/C3h/Rg9+6jk
IJZlCuypI/lVcWa8HAyJk5eQEG4UGfV/wMrDCf03URZmApJ9QCpzdz0B/0lIY7w6
3tlCwNa6LQCkaH3ltlRi9LKMV2zW67j3f7uf4GRL1/FBopTZKyE/JDv9jUt+IexU
0HUXxEdNW5UYHUD8HJziJOZpLc7TQtIUNe/y/k9m5NRrH2N2A6XOVGSbfXPkid24
YyD4x1Ryuyx5nA738U23uykKB+XERgw37CZqCxACNkh3n6uU6dbofSzXmb+o2Nz8
IXGX2Nd5BKtzA7NvZTmQtjL+mPY2PkxHYadi507PXyNp01WxdOIhihKW0ZCX76vz
m174mV9LPoddV5kYpfBP4cz7zdJKiiQpLrSBPgSPy7oU0qp8u2IPqgNKB8UEWCbR
e0UIxTVv0N/6ueo3dsT6Eqr5tk15wS0DtZbLxcqtEhnh+AwQ+TLJDFYyoY37Yb93
WglEcrDI5tApBMJqFfkYrLF2JVXpFlRN4TPB2FEDm7Ff/HLzjIJQE40cwh34LddA
K9doGjizweonPal22/LiFUwG+v+Ye9KXV3eryJvYuRmJghrlazGwgt1K2kHfrcfC
MNr2uvAGFWoFBYQBXvItPPDvY50JRTuaU6b0KKlo7G3/1ai4ZcQyy8zUEb8WmNb/
76pb0YuYQV2QR1VrcX7pDk+DGe02FZ7O+Y/HucVyGwmndzyCvenOHG1TZ+sIqeKU
8/toWtxZOO0YbxeijxdR7QU13XWEqt0S7PUoyZtcKKZmNJ+wPirIYQ8satP9C/i6
GoBN1FA/qD6+nGR0GOEbsIDG77xlU80yQe9EcjhihNNxR1Htm75HH3EHCzGNYHDy
oVi2VAtQKCxy5bBDnsO+FN8HIqpHGCyVC2DTPkJJCYn/oBs6mkQIvIlWwjCma79Z
O/uyCor/VkrsIfMyF3YCQ5j1CRJypxab8MCwSc4zC6nam6ioEYeclxuqx1X7yjRo
qrrH8If2oLEYHChNV5LNe3zXBu5LapKhaM3VqiKflGpmjzpfc9qaG/wHH9AIXVUJ
TFRtZudXi7aJZVR/ukgLS8E/vUltDOIU53W61o47pCq7tWN3Cr8enybmV9j/SqIF
GN7c0XChB/x5FhGzD4qliRJIwWECtRPUrSK9KOEr0jcYjNgakigIHoxKtyF3OgHt
rjRYCQjfPQEppKZdXTkTgOut9ZnJ0CrHKLa4/UlP+2quKwzhD2hCWWvgFHFam7GZ
eBBCL6lIlJMOvOoVbGQJ+6Xbjjiz2pcjWHhj4GsmOpGpUsh0u5TDIZzQuSpneds9
PTFK+CTQPaY+QN+tNQZ+0A3tIrVmKxeksZhxRlZwy+pfqxkAq10IKYxtX74F6Pn0
VigHHk15VfSO3GztxCie20oHb6hkkwAyFIm4r5tnzU3jkz6ivPYkBmLypDlkOzQR
/rVS+qnbAewhhyWRnN0qK33omHKhtYgZvqQQQrkiJDG8P8yzynRgrRp8jfQV0mBS
BE+Kq747wUHJBnp1RY/09w62PXvtQmN0EZGAJSjgZtGtNw2MT06YuSz+YxyBucTv
b8fvrDKgRCq9rKtGWK2RbamFuyGxR4UqRJYPhqKzORB/cw56rNq9KMds/5SGgWV8
tkGtG69JjM8usnAFngC72GrQNXJ/xRqpHIBu06vcKgD+EjDwquU4/Hq27y8ssU6t
UtsEhXd9iVmNR4aTMCq5JjyBXQ5asVACPkcLHBeG8Yt0CsH6um5S4rc6P1sys9V9
bivp3kbNc2tD9isuO0Isva1Hvz6BYWbWRUKaVW6bdvhvJb00ZhZ/8l9Hhhoe10MR
WmBxwcLn23HuHbKIYD7N6fTHztflfvlD1iCyyzYW0ljwzNlrfp08s3e0OrZ9N+8z
ifeZb5IY2xAawXG9FZTaU9i0cPMnvCS/KknzhFl9SN0EW8FH7WSC9dvYv7Db0zJg
bHA4p2guEVvjfZ2Pk6d5dD4hf/LffhCA3dRV0ju5Is0q26G9O5R7QJzD1yJdrio5
BAEGo/k0RT42iXGDs/R4mv4ok4SW3kVxDPIC5harLj29pTFnYH2Zvv9tsGsBYPHs
FGkUlD6dxqUtpVYoCHKxC0Fo3uPhV+FQMVg1ofWWCGzEv3GlKjJWcJbeDZTHYuV2
eBHTBtliA7LPoU0JLNuOShWRGZazcgI/syPkeh+JIxVuYoY2IGMV3RSLno94MeYL
EFShZPdq66uFAldEIUFtQFJY2B2mtIr4SRk9ou2wZMF8AALc3wCfco4GHlEzXXze
Y2FnJePTshwXJB9nNCBJNd/odjctzQGFk4mrm9CSA6HMkOUBjVtICUJO4wXGu/vx
FK8+K7Dnezcs+mrMffKnBp1JPkACY+sYXdCnkBMUtdd/qb+Eoh6n0SHGMUYlRIJo
7FpKUSzwXFtbq1zcRXboaTbn6GYwTwDg3B4naXaXytnDm9k+h/4pyhNoR1jt/AZV
o32Ua1zoFt7/a8LknthNHa1HPORwUip9KTUu7RqXHfhzJ7hvr0cNTTwtWivVsxe4
AHeYNVHQYRb2Tttal4AsHj/hOoVEOXvnxmFsuyVncNYd2rlfBVmkkGI4WhY8HWsR
rMUymFXHqtpMDG+O4xnblZywSXGted0TOOjZodo/Pg76kAIkRpEbu7lq98uw+mnH
TiibXEXiD89n9zo1I4ae1Hh3yY408l9Y0jKF8J0l4Hiixti8hSmqSreBB2z4q0BY
jNGUKJ4b189yU4ISaflkfxHzpZIpjf6p2ecYfjKt74rXh5o6cGJkUOJJ26KkcRxt
Q73xAXl/L6LrDqxY9T2BiCKWZH9WDqoPYnKTlyoUt0eupV6eiEBzJyFALwb5nump
FiJVVv+/sx6qdd059q6uwV83ECavAGh/HYrr1WlYjXNeP/ck0kh+ZUGUThBskjhL
TraugVzq0LzbgEH69oLROWYp3O/6h7ZNLGHw6V+3x+lYhcqtN9NDGLp5O/kaFIQP
0hsZ2diLEmRC8rNnXRIBFfabLlMPswhKyeYLgDGK6Rb96sQOL7ZBl4jOV8YbQu3X
kbdxYv+w4QrGEpgJQ8p3/G0g6lD2BCoNQjrNFa0Ezei74Qq7QnYeNh1oMqUHArpP
T6ZmizUUwLMLar0RYkiaUxzLEGV6Y1/RDXi1lgHKOZy87OZXHgZT8qjiiUAuygR4
nfPGs8tB9c8Z2oHZBjj/XiBEl/2KOJNX39E2+8z67OAg6685mIYhRV8U5Qlo4agf
AteqX4GzjKCAQuHXMC3KYHDyhOPlExKbBiIgmcH0TexOJbmU6upXTyJ95gja3RUq
cHweWweBNr8euuisbyhXAkf0J06qyMd+0W1VF2AU8NGsMBJXQj7QLqE6JnVn43Hm
f8Xm4RhbdABNsTSlT0oE7VcleScIvTf5jrkqhEFoYh7byRt5FYA0gKwS7NK1QCCt
EeR+t7yyGGic8OdCxnvmbbBMPxfIArwQdvoRp6ynQTDrhqwED+g9AF5wkwHmrhPV
IwNy3fhPpMVAXIRhb4Qig52Cq2W7z/8C67Mh91Sl1t9v7hd6HFrbXta9g3ypJ5Od
oMLK0Nsrtv1S1uIrZGQuKPadtYO0jjADEXn01ijkWhNKh6op7MLnqYSPKNk1MoDm
rVJkXygt44c0Xe1CTbOeLIhKoSK5loyqG7bM0aE2ahBjtfmH+2bR9fZnOlAjp4Wv
2OJLUDFq/QH4byc+ViGoRbElKQlJXStFrd38aOS10MJhjvl9S6Ywul2q2/yTUlRH
D6vxkR88uajOqm3LPvD4nlJb4FCAnv4DAIA1f/cxQmOBKWOZpeIouBxGP+WRJ8Yo
pW5jfldDVkeJ152ukp9y79+YtQknOHZoFeUPidchqTSbZAot5YXcTQqojPIA7DpI
h0NSRH6HjjPoR3VhbvfhlHY5MIfgFN3lE6N+zjgUKR7zmvAOyun5pOV7Pql5Thtj
yYfb+djQ+Lj2mK7eNSl5ePh87Xjje29CnorP/41W9G/drvM6kK+H9/Ap94GJIjzg
bU1KcIOA8SXFZgkvhVASBsF1CVvFZLAjwFfcauegKfZdtmC+MWk0NriX/VyfZd+b
EsyN2QO7x/CyYV/P47Lm0XnquIX0TuiyUdDBs9rRI/UyFfKyYSJXH3OVHbxUkJXe
2iz5eZcKYWAQLLYlOV8QxpHgqvy49msJjyEFE5d5PyAaeGIJVRpb8aL90EMV84Ak
XP03h0WKRSKxr6RhUm5yhHuV+0m80aSrdVH55oTqeOwbJJUHJs4xRMJQDCaQdNrB
F35qx7bjoLbqDN886VjD+OM7aDhp3rcRcdxKP/glMBUB1FvH8w2IexTtoI9xOzEw
52uN/6AGYC4NxgSU9isqhi2ZQBpJDgeJ7N0IbGjrWJ5DTalBLNpUT7ocY4tR9HHW
X26JmRM3QPN0o4SmYvkfCjRJcQRNQHbXesdT9m6U8cwMxU49eq7ZLo1Ko7i0dn/4
VWIBSA2gRNAocVy8JZFtSH6p6uACG89PJG0wQQxEW70mFq3fWl1ADt3s8UYL7Rkb
13KLjY1+lD8I8CMFRjsb0HCMAiPjCjc14CcPMHxWp++cmpMro+DhQDLCP/Ia7NQp
y4R9hx4JW9Myxi2TnuayYgh1Dm1xfElcc1VAlCNeawcYdTHIfVUS7IUVSS9Q3SKc
T6ahKtUl5BgdIECTBFErcA0BvDnFaN3+nc6VOcf4RK0BrYjkhgo/SGSd3U5DVABb
yMFKOVCz+ifuM0TPbfHXBNXlL0HWLbYmJANcxoTeaWEfAAzIsxa0n4eTr3e/kgkk
n8lxRJZMbRMufW9RJ/b27TwgXpF5bXM5I4yBm/h+gxflF/iftSxWdDO2lANb2h7E
0IaH/witZAINT83X3lnF0m6qUyKc9jXse7t1h7N2Ea63tiZehAWcnzBwI8e27sox
NaWm+ZTuUwgxo3sThc9yozFUTbB2yrGBvSwg0fI8X9R5+5hrosMiXlOxal3QNgvr
hAkshHBFi2JyxIDPWhF0hp8ZfFDkEvL8R1OpFgPA72+Ecqxzsy9teuOHlaDsPhVw
LaRxUB8qCqX6RgJJ38meaeKNXMj5/UEn5ge7pUFlTmd2LyWtyPnV3kYj8A/ZwSPG
VuXE2mEUhK9i4yjbO4WIohwR7NxOgLkFgROJmo61oMj6rieRguVljbvxiQkojPDM
HcVAmL8c5KQT1xhu8DJY4AhEB/ZvlOGLe8+5GaNAiJRpxBdUGYYSDCBqxu/cEQsq
4DIBDqL/lgbh/R0h8ASOnCRy39VmbieCFccvqHIYWwo9FDzy3uoxh/7urJb1oKr+
FGAVAc6kuCiRCihr9enBOi9MySRKEZ/6K0gC6KuEHg7Ylj0uLpN3cVxtAZb47GTE
OgRJOasSNZzGB9BJwozLqthWwWSEbtlLhQdM+5MhiXDl4JbAc1jzBP8klIRLmiOR
SMcZUsQ0TQx9eH7Xf/frB1TiLZFse4uUbdEuvO4bWxIAvzkgtuY18M1yC4aUKKKS
7p4chIqpKCTjd4qiXClxUUa2OJLiqA56f2WVYRqlSR5s+nLWicezQyRmsQeX48TC
sd1BpfEOboPNFxmMLKyejHLNZ/NyhfDd+JoFBCoMvtIP67wXuHrouRoLh5/Y+4VO
HGtSoUXkBPVqXPocfTFIwIxPQr5z9jhYBXF40aizn37OOb7oNpEkIqHLWM3O+2qN
fPBys/U59BCiadjHwj2HjyJxrCa8cjtyEma3PnBrq6TGOEKBzYqegLEVSLiGmopH
aydFqYnoKPTlw8UsBdBnjoKjlIaSJPloLUxlcyt3yC8lLxzXb/ZCXjEIn60rnl2A
Z+PJXkRhZTNvG43lI8eBl8O+UIJNUhDXfIaFwNspTyveSyG/3E2nSfrCaDVRYyZn
ZR8Va091/3QpQFKgECPI6OPlQB4PVadXEE/K0I8L/+08CWj3oTaI2OyuX9Usqp74
CQYOSTbk3e0hgs0c2gs6fcQJ3+DS/mou8z6vy4fQyFiRCw6QbZe/OOlCgsQianeB
QMnhx6xkaH/LVwVeTUB5rS2JT2mJ+UFgTt5ZAWIDcjoV0PQRjBAck9ZkfiLLjYKf
zOB0xkwQy5/56yIGAuKpl8B/hafo93rlCMUyewch5F/yhSAxLyAN7COdjPqXvRAa
ScA8Ag7nIpQ1e1Kga+Ue43wxYDijDkCL4eUu0zY+jjAJaCtgz9nWfG/Jd3VmX3dx
ohiOWTdKtqqvqUJbqSN8oTekBX5pwfOQmTnaoIgDldunXKcSGcC/sSNn/3vuqXoX
k28bss5dDdW1KWOfVflG0ZiDwy4jldQUvGeBPMmkzyjsqCEwurmuBx3XoIsbN7cY
uZqQuX0JeehoLV4OUHpiIS/rfKzRS9RKyVjy7oQRC630PH8kxx6px7iEGOEu/iA0
olKXKjQcl1Q5nGRzv7UoT8ra3fazOZHxjarNYziFXdMqbyzh74n8mK22d4WU//yx
dhaCqk7Op/+Oh2623SwMTHn5QaSlIAaNYyMnyO2+yYh/6sNiYXij8fyUi81eY3ul
QPabNBbFRRHO0wh2xbjqNZZlpBFL+4cQs1YKlCmtBquaOHHBrYz8OrnyvM9MxOka
bxY2V7a3g+6O2Fp2NfkTeRXt6Za6fjGUCE8DA5Ztb1G7FHCErTwQOF/2ztaKnHAj
pzFHcltxCIf2hZo4aNzbN4YfVQllWot64wJTGG4d+KX6FYuWCie+Gbi8yhJC1IWt
51ZO80hI7hn/yr/8aAkBUbcB9iTMKskPha1Ugl7DsFKcoweUAvQVul50FLicE/9X
bps7Hf6xTWzVGsW0rjP7XAtQx3a6h9KocwOeF5QB+gqa+/rsdtqBrDjjtTP10vW6
dmiBLslhElIbu9CrzR+29CMDBZhFDbfkuuCEtteZDGD5pfNd+wtp31+Av0lrgb6q
QqZcdMpXsIRgER8sxJCREhOPepOWyodfW58qyXxugV+boUmfS8iqrqkstB4KeMw1
kz3m5T8m8+o+HvwziNSqGkFzCQVdMwPOO2SS58cHuv4BWBlatv15BCc9NMBG/s/R
Vf1A3SZF+Ze9C5Rr0Q8igGX427LuemhfLtgJHxBwA5ZaqmtrRli9ZZ0sGkDT7UmS
vnM2l6O4FQ7jxtvfmF+5CswBEwNvHglkD0DOVFzDQKTjhxXXVpShyBKHhDRei+q9
Od+9yirAP3r64MFYqlKVTCREMcISSdU/UVNhHRFH7vtULqFZfctyf33Sby3D49Lg
3lTPK0nmBa2TmrwF6YUA63tSwkKF+lZcm/3XysaUw9aiYKp5XchNungaVr1joft7
RqpV0b5rCHUzaiUau6Jt1PWamZceZW8CEtt6u2n4m0+I67UUyOu2L5ka/8wo1AtI
qA9YzMRnCDA/O2DE1W78Sl5T5taQSz3+qxskpyEZja8jga9RQdZ012QII46FNAtM
t6f9mYTVlfwBVk5k584u6ZpQQkTYKLnQMC7ERyKARCsZ7FYYLDO+XvHiXtK4xfaP
iYp9ndooUF6xd1Vu5WZHkMYnF1KQU5MfOb9K4XfU/fC0lVJAZmaey2J3SyfG9S1Y
DtNBSW6s32CLFZztOsni0PcIaYrDqXW92WAKWgEedwmCYbpJJVkuNSsXvJsaPfxq
Cx0MLmoops5fVHVXay9wwbukrNK6JT4DXE6rqnPJl3t3ZKmnQFdedr2nJGu7AGdt
p0f1Qvs7OEeT3Anoi0UBhul3JG/iPyFALmSw45T8uCeP3YklCb53x+qezrUIZrdC
yV/epUbc15fyEWH3gaSXdzngiUABAb6+lHvs3UCn473iwDBe8Y0gGoaeH/LuqOZs
VsACadt0sjciNO12rIpwkHKsKzj0pb8Vqv/1QqpyL9yJ4YUns1TBVIv8n/xfZvFW
xayvnGFpOg4qcg755DaXb1IrxnGB52TegApKxh5icSWYFOIgXCdioiQIf9OYwTr4
ZzUPq53PG1TtHDmmpTHvYXeV4DtSf0j0fzJTZDMHClFDKn6CH+xdNVJYv9kYBl7n
OwdIpHplUFU7LpxoQXXyGUnegYI/q8ya/k0riV5ehC2NMg89ZYHAmZE/mJWRMFYJ
X7hbhAz3tLzgllxkXpeg9gajwXSUOviST4NntpFfMC5axRpS4W/MKmOsZYwOstaR
OMDBThV5XS+8AjuccE6vuNbu/TcN4eAHJcMrBIwiQ1PEr+Fm8TueqYm6HhDMMdso
f5zhCLcokikDo573wav4AqlXbH4nP2QsbdRRmr3bDIruy3FSMeIgDJx//Zpnci0I
QoVqrGW7d1rlKuyc3KGiNcmbfs1pYqGpKRuZrcP5Jmf84k9VGXN8HxJb9BhNMrdP
8G6sjAoNYYg1xuaxGcZBwUjXkfvzkTq2T8X0mz6qc3yP2ud1IF23WWuIXpWBZ7ud
rHWysXsbN4HCcATskJJGWY52S78NhBmkodPIph37kLeM/iRTIgv7U4j6KM++iFXA
URH9lpxdFZynw1UElCxMQOhy3/NeOPzGid/ZIEsLuy9jc2KqWgPR18M4i6qGeB7T
s7e5UpAhSC2dDNb2jdqFIpZ2XYZy5kiaj56PN8k+uk9Es4QHd+l5CKD9NwXjPXPa
zMhYVt5pWKsc06HGlG6B/CZDK/D8g+HZ7tz+yYgIZpdnPsS95t07kYCVOBAlld2z
6Vyw/45UaqQ1OeFxdhEsZj+lZgYBoCMVWA4PgSEuESE5MJYfj+fpFdHbispk7hBn
y6hVq0yv9Uex6TAwMxdW8XrhSZMlJTn/04ohBa7EbBZxjwsqzqKfcpGZhUjT7RjY
gX3whenglGxEiWav5CGzaYPBehE5vmXVkELaf6i2HcWdODnQbEaZTAYuRk7y84p5
vD3eZ/tURsSCFYPoJR9QsBg1kRFUDJvdq77UEH5A1TugRu08snQIvL6KZSSAQAhg
HoVbX2+MBEYEuQYKLsGQI1xQ4/Zx8mqcSSFzK8VYfKX0qE/8nANJPOtKr5ELJyer
kMOw4ee3l4tsT7CeSZKUlB2gk2cfgGB4FWxKvIYAg5PUsUYWLtJFGmxV9XQ4C1i1
Q3y+0RhiA1Bjh/87g+s+TSiW5Jzfap5eyzRQB2sBJSLwv6Zmvlm8u6jo6rxO15Gg
AIFOe268xpeiH6bt3SGdFEblHCzDfjFbY8ZgSGBwrIwl85o8b8nmYV25xZNgqT4U
M5z1SwmJ5J5/kTBCu0+u3A5dszcpOt0/1hpFFVofyj721YP6NF+QI3efOHILAN/F
v92jEf/kkKwHKDKLIWVq/6NdmYVlrWKoiZo1BogIn2IpHNqN87pjx+6lV48yAt4O
tpip+dyrrA5EeNA0ydAVt9ZldcqsSIo4ZwKrz7hE8OQvYkfAqAYW4bSvh9P6HoW5
Ka+ssAAMpHfbzs3EeA73UsFIJIYWDgm0x+9k3p+hLUDceUbe/mZWuTqbqWMCZMkL
Rhuonb7Baqdk3lRgp8MHaiftimP71fxvsymt+L4S+rwXHX69SLyc8TlI1AWtY8Ux
/Jx86edSMFYMHUrER7RGvS2DbooG73m9ogd+ElLx1EkrnelsHncLXp44ueqM02SF
noB0zdG6Um9Q3Eh7reu8G2723hEpvgNzqxMuPQLFig0oEce/DCwA4v2pBQl4AcRG
Jr+OtfebjGhSYDvX9hdgjG8N784zyjMIrS++5TKR1zxERgDVl+iuIpT8ofcBfURU
2jZZYvPwOjrLRlrnaJ3Zi8HR9ql/DiXgdO/FYAA8AW+JudnHes2npOfUTLUQqeGU
xQ8GyaPM93b3uOh6uY4Kl6cojCj/NdCYLKNe5ZD8xW++B7p9YMU8XCaFMjzwViMO
CPKZ0YKYlvMkCbYQ+nZGCgnUQD1LFlnhEHCHpeIz4smJIzC9tGo+Hrv8m8rIjqyL
FQ/HrB5dJ8MO2Ht/2sIhjSAjgOKjOfMWYl7xxSaZyxpYcBHAb1fJT2ZZXA4KLd1J
y/0AAtr9+S6FCoTrjevVRtZxJN4ZroR3P64Zscwv/125RB+Ak5YYMOQjjh9X4+LK
7a/Hz7kZ65j1vQni0K/s+ogKJDZwWIC1RHI07+LaU+s2D3SpjFXqXADwepPGfMnc
OfLye7EgyeJkLAbD/OIlEpFSxqScRdkzQcxspQQMJCQ8SUz6kQYy94zTCnOlvUFF
DkZmzl/1AT+BLaABYkPIhkHhky0AtIohwM6yLdJZli47MWPPJmBAFQnPZm8JmiKX
g4y4y2IfyLP9JwTm9SoGQyxHqJ9k+VrSr8Fmr2tpcmmLKPzkJrZZx7+t+Q9CcZXP
t6bA7bXs5W3Xr2hxCPZN42EztnDShOYud8//B8t8s6zAW0UyZm5WeRoFWxahNh19
8X23S9sp+rsbISvMi70hTlGLHDgl9qafCkQkYwO7VojnjIkOj62VjW8Wq4yMwHn6
8/k1BNcY9mmEV8EtdiD7KA7U/VYvnGn5QwTgEf5G+sSEzIxxU6nLFYDHFjOQ2bGM
r+TeZ82NuH2pArnDnbQRF0LPeLgTS58lYcvR0ZyuN1A4cKxx2hlI95I5imF0jNdr
uLEqWkIVHFjI3aj/XqghT2SCbe0n7WePlNsU3H8oAqvZJcuKDD1tvibJrtirF4zL
n5OWsRUATgZ0VKccoLN1LnAL5iQJsLugXQLA/Xj/oJLIiuMQRzPK17mgpe/kA0TP
qGkhqJPTHa/TXVo5Zk6Smij8qqPfYx+/RQykWpuDTGf6rsRM+GfEDEfDWNZBYv6W
6I4sv5YXaT0AS5ApKsxo4hCyqKqjMhCjMz9kahQttaCj/sW5DT4tNCqG92/XooPn
PFvkfOmsYRsWsM6i81YFe3Gwh09qU9/owJzBZbD367+EUoc3y51JRngVrikkxP9P
GsR8oSazc1FiaMJD3RPskODcFkOya43o7IGd0L691TPYdx1830yWuTCXaZZd+RJc
V4xHWwtBT1LasLYUS0T6tZXSC4NMGzXNWIBE5zO7ba1ZVJR/gL81TSTB3qV6QRL5
eiCkq7RM89Q5ZNJbDy8WnWePouL0c7kPfrb+A4OSLdFdfdje7AH8QpN4pvFOQrEV
iH4UYKEH/PUf9fPBU1YO1i0KvS6scHtBLRks0NVDm4Tz3nXDX1GCz+i2nsLFjGDC
l3X2ANk5UpWn46QIi6CPZCZHyrU0QERE0+01Vl1poxlGRsvwjhf60BAeVeZPw7O4
hTng1KZXnwqUAQ4xk9wYjUyhPxHgHcCzJ3PzzFuiQJGNci6CRQAI4KLG20+HgWu+
8R0IRRjJq60aAm+7wiTv5DCuFeuKiNl3oJ37xsU6ZChPXhrvH0GnYwPUgxR3ZRRT
y5iNuSjHcZMzqb6T6qeEmvZIpdQSbN8jBh3WBPChJzVj9ZVhv0A/Xk2GeA7elIJT
IL04mvo0nHh3j8R/cn38ygwz6/hF0gK3jWp0OpbvEXpaTY+thZCD7hwUwlg3lzjr
shPMBPv6hwHWZumTodChZKafGqw8hKvfWV0ZmP6Uazs/7qwvDPBVTbQ1BawbhgfW
/HXE+VwfwLEtuMMMrMKPCw6OHA5dV8xLQM1g7eZuz8KhUsyRut852TFubpxCXUKk
nGP8eCaXTthoiuH0RboRGnk8s15zuu5FZLlWQSAR5cSqHd0vnf/MFB7km/czNmZS
uvcE82dN4moJX/sz6poyBi2007qEnUdYj1VbLlMeM3H9MvpGwAeGLaS8l1jQmiop
cWz8WscHy45SfRKNlLgXbBYIS+FZIWCXHBp5Hi6TySKgae1RedWdVa3zJRT+BemP
3gxZQFeNilqWipiQWcXjBorTZ73cHdzTC2xVHLzKZfKopxsRIMiuLHKqO35BkrEE
s8B7qmAi3Wp4E34iHru3Tb6piK33LEi1d5+cLU4nRs0/mRWY+BWXaYwgBfZVdVE8
C27fHgYG3jPdtZCLapWT/doanWMFb6Blwa3W13siLEGNZF/+Oz70dckRu0GLee4k
0zpFA5GZOd+lq3q9/4y74h1JTlD3nJEZ/NwJ3PXCZTykrvf/rpOv0OYDCkAQmGR0
Tyr0hZXukCCM1x5Lfy4uACRb2pqqTPzWf/zfASdundzn7UXUK3lPVdabNxPg0/1I
Z/d9oaoiz1yiDAzW1jw1RGOlLb6rAZD7gygDq+OkasaGfqt+bHx+eBrDz/VWFvZi
vodKkJdQb59/oGvKMSKnRT21WqNDeEA8hE9uuOD6K49rMsxykPvBeNSD8ubhd3WQ
tVSlHd2ExQn90B/fAkxgF8MzXIYlgHkC3xxEgyVdUl+3sHAbZc59M8g2mttblldn
2ddOzpZUH7cpEUdp9FOjgoy/PFiJpUDJkQoshV87CRxsoM0sa/4Ra3oftRd2A3dE
LU9Om4SS+DnSTHdP3bK+RXFJmBOO4f5cU/7h2GS1vHF81s5BVf9hpUVA7ssOUU17
ZetX1fbLMnaqTqZQ0HYUA4T1h3VCMqYZVtdtSQW0d3FKmT6PjuIe1NQUE1hfotM8
cD/0QEghr8VIeReV3ehV04vOIXLwkax4q1Didm0nf+T/udFRUzD8x9FRI6C3OOjP
z+e9N7s4hBCGJpSoiApUUOyTKjiZY3xwFh/BdhiWT6iev88WyUiIPg8cw1rL1osI
n7hNFSVhUd/luKBhELM5aPiDfLhUabw0qIk4hmEZ8mJsJXDbR2tGjUrRlsdeQJAI
PhmS6ePQVmRXesnvgoO4mXR3B5JIXtIMqfxmUuwyD6wNYUka/TbJZFLiyeM7GOVn
a/EG6gTOo8z+JbA5juWD41JXUBnq+8oi54lYNrDLVrW/8DCG82/kphWqDMbKaU8F
qHNIwz2WDPEE82y6NgQ4RMG45J04Ej8KFW3dpbe5uoIa43F+Qudk+TA4qcpEooxA
eth486fQCIoMrBBhu2Js430+XezHsaekIE6tXA/bxOcpXk3iBMXfPKGR6NMxfzlF
y+7YarPS2Qd4Zq19MiYSrT/dDa86v+PaW4Cls/PjpesgOlORwMdu+ZsAxovOP/Va
TbM1DUFEKMBmozp5I8HR0d+C8kzjEnnL68Eg70bnoKtgL/5d2JoagbcoBsxDRCGF
Z+yMTwn9xhfdiyk3aFwHo91Qtu63bhch/niHY514zTxMNPIvsErwAwDDAjVc1JST
henFIZU584ZChXCoVwygXAL+jn7eHbEiay1zuDQPY2BwR9+3/LlekS4D7fA9rCZ0
/brfPC/t9puHsxfyxxIvDZw6k7EEMttY6UE4YvQqp9TLHWg/BbrezZmM+n26rZQ/
/O3arjipkBwYpiB078d/PaAZh9tqZOVcm31zU8zjzjJHacUpVosrow902keyeDhI
RnTr+yENbwQhrs/RH/4/BrvIVaH5ILVaZh8dIOxkjiFd9fQJi2+rl/IGf+0u11jC
MX84t12FLhmCyO92qAY64AWAY+5K826lf7FpROJMtHuVIQskZFXTFMexAm2Wr3B+
2vnH/puRV19Acyov+GP4k18Vq6sT2MF3lxnEr4+zJx4R/AZT/kjewKP5oy4JFmlH
JgS4+XJ/A5WNhsG6ewtOSUnJlQcNsHxn927T5v3hKPJMMomIdxhn573RFp9iRLGQ
X58ta0D0b/jZCj3IkKfNn0+84JC1/8O9vBKiA3EFLbtpyqe77MimNshzF+BxpDDw
pC7r021Ek1CnMeKyuN4oRaeuBifmeKSmWuZPIvyDETNqnmdAoRVGPsD15zVyJV6w
CGurS5jGRuiYpZmZ+RxfX3Dy1JEHmEpT3FErl/vslxlupWMyLIESCK7eYrehkmLD
FPzPfFlUutPD5V3tRvghzCN93DZUUu7fGm8LomIT7RFLnUjrC04qcSjUImNgGa0c
icS6wfXgDW1nHew0U2hvoq2zOrPwXFKTfds70ev/U0w8G9fDNAfZJznAnFZZIn6J
IqGbR5vgW39KZwb/NjZOIJ9UoHBW74ks86siO6Zm89u5vvdFDv4pT1hKvErBmMnA
YAZI7jyJJmLgz/SCiDqOT6D0qNSxHs44acXlB7mIir4i9lF22LJIKMdemkm8y62Q
oA46Y1k6CLelnCs0EmGP21eO3BTNZrjGhbbvjLqqw9v/rVfC2IXHAGDVLGgt9qZw
NBAWyS4kri8FzuD7ImWaOUPbNBwOmoqeWXs6fYeFNaR5YIT/+kt2QE2F4ACJ3OYT
E9xZ1wmBYarXkoNy1zHT5b2mJx9J2Z7DwjK+vWn8jHvAi4xyq9EGrCRutZLiIVGt
1jynfyWGUgsebOba0sDuw8wZ+VYEbGWDS2/ZqOf1t41fjnEAraohvLPNu0aDDA7V
SaKLWwtHmyMu6G3ocZ4fONlOPZeRNjnEhr4uk3vTKtYm/p2WdMGrlRdrjG2RT/RG
kSPCozeJc2/ZIGHNTA1ouu/W8GQE1wNX1QcyNP8vJKZUmCTIrj5UjaJ6YA7gE3X4
n5GRDDJzw6ZF8ck6PuDxRAm3DodPRAR/wFS0/rIsoxIeFwu0G/MTO3ARpJNr8POq
BINKP+8YzAsnCC41OAVvHwpjNDsY4JYmWTuHbvjH9mjUegVy5lcCwqpAY66p7vm6
NlqbTyoPfUWEJfMo90Zej1FSVxCyGOuVeprxnDrGzCODwFsf0usyKOQ/mtv2lONj
W5+AFBoKpZerhpoh26fdhWACHrGHMdlyN+Ya4N0UhdCEYAGEZPb13g5jgszhYNOu
Q4BYLn6lsCI8T3HEfh+V56lmYCaigGz9VyG0vO6911Lz2zoNR2UdOCepVuT/VbrH
W+WV/BJYRdxTyBw3R2k/6XswawuuyP5f0JRbSLvxkDjsnggwwwWGD0jz8lEPD4XL
S4Ve0WQ1JX5VMHpNimD29JcAnR1lzjCh+pd46TUbHyI+3A3JdLERpPNLYxRq0qcZ
fWYTF77nrE7Edhv2SqDAy9EkKeOP4kwsqAJODAhZ6hSMRFJNNav7YftseyrCQYH2
PoFmSPLCyz6kwe5AuTyUs1cGwrFvGeeJa6g6icpVYIOZfTE1oo8qI81sZtdulxeQ
WQobWaRjSEn2jMyIe53N5iYtpvppohFcCBzTEqZ6nZ9yksnshRZmwiLS+6AqsIzx
GJgCwwpRYuzpMUv3sUEf2g5VB0Zx/ohrdOkEm4MAdzQDk4yDJEl8SE/chtaLRfJd
WOJEgkIPyz7bORrjAITMb9yJsaYputx2aSj99OPn4qZ3qrkEgtTtGoa412dkJ+XH
gdPMTogHfsixuXznKufOoh+9aAiOedGmzqog0NH/0yv0e4B+R+Swb9OkYJLBDkX6
+nMeadVlEo8wVo/jDApkieQvhcKD2sgQJz1U9k8lhNr6/JOwUk56ywchf++gcPxl
1rGjxqU4aPELUgbV0tW6aoRb0+IesxvmfwsMKtK8cLlPHPt8H7ltwRhgBJDy8gUr
MCXXFvGx7UOwhQIdfXMvQOdN739DtwGJnKDlymZB/XtKJXEYVEsaSeVDzQK4jeJS
MmmTtiqe6p4U4a6I3Q8rTcMf2GeR4+6Od0FVM8cxcO4vpD1SLck3q3oHEZzlARs1
/FNIr5zJ/Ut8L0NfzLd8UG3qaiAyMKkACLD4+vEHu7Wkd8gePzlMd6Dg7mzOuXqM
UfRdeLGyp8nnnLNY8XIZDOYfZ52I+Esewf/J9UCsDiiQrqK2fFvmrchI2PsbsEco
EnDXrBku2XbUDvZRvTd3Iko+h9l/1sseU+HLckUxRsjDrZeS/T1JR9+o61lD64L+
DcW1SwZqOfke21yO40p2+K1ghA9oeEXQA3Wu+u/9m1odkI29qoU4vIOZgJgap6OB
phNWDI0Xu6fBXgZ4spq4kgM+Rd9cvIU/AMVCApIUTAXpK2AC3ZfhegxjvZ1BI+jA
xIOiY9m31xxrR5quy+KZQ01uDpc5YnWxPTp/wwLM/UBp+PNm44d3ZcoilzFhcS0w
ysh5VH8FkO9zV6bOh9tFUn02Nbrjp/H7yCJopKo012Nag7cv88b6fFOA6JKrJtgz
Bm/RFx3i/uox3YNha1jlJuZaitRcywXmi0g8AhnOw29x9fT1YZD/F8tfIQwa4LVZ
pwgZa3oB2xIGk8I3tL2Kt3QTh6aBs6+v6do670tXFXuqQ2ZUkOHNf0bRF5kn9YKO
jyneV78zJGmSK5u+Vr1uy348DvvFc1TT6ALTOJIri7QRky15CIPbqx5fGufDm01i
ogIJVejiIqBhlMX9x05EW3XCwt1R8GZpzKGYCZOs6GQun8SHyTscsefAddH+hzaV
KJfwGDg/7zgLD7suvpI9Y1wo7dF5AVVGeIBp5MUgl0EpfeaguouhXEiRyNsiQ10I
mseghR22ri7uhEz2qJy6I+IsXuP98E/hMq+BAQZHOzJGoFrzVsPgFFM+ywzkDz+U
93FAgjN8XioYi8wOgk+bYNsUHv0GyZPhoGo8ImMdWGLivkfbDTTzEtllDLB4RNpG
GvPWsBvhjEr5OwpGkjVTRRtqcXiGg7ReUleq1masrFgHKCUQWj9fsrDxXUfivUVW
VAetq2tPyZVs+hHnOvWuXPKaUdxc2K4VbAe3gKyM8mJBVoR7YkJXq0EvsmOiEF7s
kKyzSmoe+Nw/XHaRcRdzXDcCPC9NhDOMwGhPgaYZrwPcRbSSrUcw+tm1stGgxD/a
CpEixlJh1RCvYN28pQ5FlnxMX2Lx3wmEAkvz5N7E5yakAcLEoEOAYsrt5Em3XTJ4
RbwCF0ED3rt1hQQSHiscp5ujcJFFdvDGDfKRuMXWR2diKWxAMh+Xt0ki0ZrL2jTz
zn+WVcwNYZFvGZni8ZkoLf+sgoGxfhMSJvOpBx43R3UzpKTIF8DyJx2ysj4aNMp2
j2WVjJzBxRYhI12FlHqUMBdFWvEcgxM1Y9JYLNrOWWT/GjT+Pejq3dItLBzOTopU
x9FM+OyB/InCtltLnTNsH/srg9HTNciI/y9DghtrbXPpZ/o+SFB4eK+TPBI+JWmv
4dtGxY9i3DO8LyMvu8m8qAe0tJmeDzhG210jUQOK7XH6Xqnwqpdo5dt9LfraDGdd
VVPPppqvClKdjwcJhMp7RmG9H7oQhmFyRKmdHd2F/k6+YvXiHULqHF5gohHzgd8W
l1OuCfwpqdJ6vKH9G7x9ALa3K6RJ0irtDWLu4nLsJpmgMnnfXJibstMeXGc0kPhw
LMv6VNLd0CeFHsCXDsJbj0BY0uS9JDIUT6B49BNuxpXa6yqWTQFgu0S/vget5jiM
f26MGe/ykNTrfmrOEb+xJUs9Xzl2c/Lkw2Th3KqmwjifgPJ4Ov6Lpe24d7kO+CuO
SQaPtzz9y29t+HjOeF0HPUA0tXHN4ozSdNq0uXjms14ZMs6op7/uarToOga8auC9
lfHbz36V39UKZOyV2lf3RlQvAxi9u6j+sjNwe4MstxyBRHA32ErJ6qj4Udb/mTYf
PFf3WEkt297yqF2yMPropQ==
`pragma protect end_protected
