// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FtuTk2RseJ4RSBJ04v+LSV+M45SmipQ//LRsxY9IKZgp9bIjSVPUpijJ0Ccjzhkg
6Q55jDnQMl6PMXRggxMT0yImNDz0NjMq5tZytFkn5sL0tEJ0wj76BLRiZk1NSBlN
+9ZPb2uFaCG6rYRsMkOhB+0M8UWv6vTnj0oEVzggHT4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4272)
lmFW/WOgLjoiHaJtZsFlJRwQzxLC4NXXOGmGzQluoyiaZbUo/1TH2VFBJ8F5YcAw
h3xfK/WEwaIzxq3/2IG6OCdvXOaJimaeGibzzMLS5gpgMIV9nuHebZ/wdeoxvl45
3Xl+wkMRkQCxByFCyCP8I/bRsCK6ivB9iwxRrOHmY8Jo/bSxfRFwQIHl+6kCy8vx
QTOVLhRy8voPNRYgPdfUT457/ulv0H4g3gmn5LQ9m/tNt84Izl7PM3dVDwZcy6CX
PVAXEpQ3kwBxcJ5j6221wepYRqeL9Ifv6lNTgqg967hEH3dgXoTT3MPPmpysA8Cy
FP7f02GRSolF2i38OTUqwTS1Qrb70nZCxrnbVT7YKfMX8l+BL9nTQb0N+NaxPeeN
+9v3dx6TOPd+R39a6h0brN2MrjRGbasgcZ7wrsDoHVMRis1X8kF+KgI5oso/5fcS
WgByco/LBASpQXXCl1ZGRHcmDTb11amSuvH6sL9oeb1/49fUFTXTxMpMGj+UNkDP
T7pPeP3RUdCTQmH43jhGYvQKq521zejMndBFbmyXlflrTQPgaTnX+sRHkSWYcL01
Be2VFepSbUn6K07qQyMbZHJXuEJ4F1mFDQ+/CLB0FwattTCG9tHjEDhZTEvw3pAH
D1JbbsMuU+V0D3fKtN3RsFhcO/WMr6Otm8OwQhB+QzB04298zGSXdBnRtAEOfhXr
pFA9x8AizNnqP7QK1CbZ4GDsJxqmK+fDOXllWx2GGIv1niS61ciMFCOA3HFV2fyE
G2q7JV1q7r7SYuT2pz9z3rltSCojPJMrvpmaclKs6JLnDLzcfMEAq4fNb/74F10S
bnufhbMM5ELC+bs8ot+qBiQYPhOLSeSmv179XEqw7AHaSqWdXKfszmJZvOUZr2z9
Hsf14JQ0HFOzHn6XRFMdUCqu9AqQWDQydGwV38DkYMXJ2bh5JZR0cmCzHqDAEQWy
ETutYVGNY6v++6GpFNGbZgDOQVQhz3UZaz36kCCy3fHvUFrHnCSKnyGky+fSAqon
SUUsRNl4ktkYKlp4l5ds/EhCc5OSLNIlwe3NMLaANngNMnCruwAjMIWXTCFYQBBk
7l5+D1n4MnuH9ogCyUQQS1dUruA9L4XLo5e/fc0ELXBTD2yVxM3K3JclzM+hReto
oMsuwveP5j3D5WJ+BZ8UxQMcf3B8Kpbd02RpBPZCkywPCnUDeuj6SlArJjYqaJCI
e2ZtvCJeE7pjAywxToWQBI4CkC8uoaOCjMSELk09VzDWRbEaJI093qk6PjWlWyP2
qbizEtSCVKnnInzXE5PPc9erbGVhsCcbho4gyd2XEjySmJ0zJHIxk0TrdX4o2Hon
YAlzUJdi8/NHEfsfSA9rIExH2Q5FpofzkOGRRt+JQNCIyBAjw2wp/GBOMySeQJ2C
/+z8oNKl7jEqVx1Cb4IL0lNRTn6qlIFNw2rhl9x4RqCIK6RBKZI3lT8wRRO6pUz6
v+fzhh2RNui7OMkV/VjkjkbqSQ4Q7XOfF2TAr/7aDSJeDtvNON1m7v9hLVu5AILh
9ooMVr6tpqfcn4WFMqivmXd7bATGkAXU65hiUIM1WbHsN/5QUmR/P8xN04czM+ot
Xa/wjcdF8g+CzDqBWDJiPySZFPWtlmm2N2F5vAvavpC5UatjotAsfOpr3x/rWgi5
Wyc0mSrcINkwXJWvyhOBNRAR4XiSMiwpFzwt4cA1xPqEVWayL+bDDni/E82t9Z9q
3gCp7xbifUZEKE7LTNIwct/7i+ZBZrOFoUS2JKQa7FmWXlL+dHfiWILTD11JchCI
POpM1Bz+qmETs2d/tXf+8+GTjTplKIjncdnmvJkdLoFOF+PmogAKZgsYxRgm6wlX
U8MHAeNcCcuq8MeudFhlslLsUSAZgo92/atkOSLS8QMrYRtqapvFAsysfI/ziu9x
sqq5IsbTA/f+JijWmLttWs1EKF7Yck0nmPFmKpBqSKJLbhbNYaHnPQR/WRhSkro6
IZ5KWR9xphTZudUw1wUFfdbgKMssD8hWgSsQQmpUBrsC0MrUnwMdsBMwKLXzByfX
2yJjkguSmCaZfoOAWI4or/5vkbOxByP6URXORYGR+7H/TdQWAJ9tgxc+ELVPa1t+
vx+A8CUG7muPC/j0ZrGD9KUMHyQOrYwvvA/VIfEW/ccCua4+Al/XYHS3MRAAnLr7
Bla2+Sdg6RTbkGGAgfy97CjDt4iG/NVIg1X6IYaQoltXhi1xxSoc+rY/2WANH11+
pmvs8iiF0MlmyNt0srVPb6q039ho3ViFyL0+ItDCUEi4jZGfiY2AAiuAyyRE/L63
A0FcXjPjBECnCetiTkmu7RK2IGZ16AIJt8BqPOiQWJ1VTZWELMY9A7MbwXX7Y1JV
YIijQdoV8yv8lhdoqVZB4fwiWseS69mzDnMJ34dcjF/7PVoCQC+plGEZxTxSRL7J
JKefooXODZtSNXbNIuK4Go2tDOjXJAeJp6idFRjOjKe13x+A/ANeZxhKXQQyfPm8
zHNS7cmDRctFbYJc4Z/abyrlnybo3gQEp12IK+onGxtL/EwT8lj83xa9pn/8UQZT
/6rj+j6HMDkf6EaByoAueegy9duP2tvYvgfJ92NVqpy3fLeXWs0aI18nC9RKNFjo
6ZgoNpeTbuPSKc2TNqVttNs0Q0fG0yQKpXbj6ZHQtKnIq4u7Bqo2izcYWID/R9xZ
W2Tk8JgFu5ZpOn/csQCQT5AgvQh/wCLpArPbq9JpmiOOfaxII78yX5Nzm8ixRwdj
erBYf2NPN9H2+yQOWEsomfqnT39Hrx/W346haBq6f61p+ugHQDW342VqnaDQRYMe
q0eG4i6X/JVu9ZS028/BNYSyTkFV6Fa6T9OI88OOKSwlh/OHHJCmiJP3xc8MwhrZ
B1pzeRHpt1l1MMWwXXtgds0NL50+ZyivKtzM9avhH9SH0/JlPgdfdFAGXjvNZ4vr
Q3rMUePbj5rujenK8QrAENYtvL3wViubkVlLMMGWw3rD5mG4+2PuA7c1Mzpi7uip
MatASsERR7Yp8vl+wwJ5cmFjHFeEjJw2EP4kh7GAr/gfO3rW8EYzojxZgz7rkJEh
wMRzpXBf5xH9QrpNK4pzPM6zF7ZlpMW0t2w9U+ecXATCwXyXtY9c5ImKLVqB+Exs
IABpKvcZey2Z/Ey6ouh2kCBE6Tz4VJghlZktsSmC7bgvcxFBvTt9VoUC4YSsPBH7
9KP/3ZbPbiA1riSO+H/q1cTFy/vGu0aSAQa1QlMco+ta0ST9N8Zo6mqPhenz6zOD
YsHWo2NmcQHbAwwxSqY4u4ImdPn2MVieLWSZvNW+shPt0P7iSgudGyCG1wP+WuCK
ys4qT/c9c6fQ8x6H6x3mpKBvUjJDNP7Nu/HGu1lVt9+dcs6Ckyfy/OTVus/jY3J9
UMYvqjRW/TCAWvu4LzjW4hitcAlhDo5yanxdegqWri8GWLipfxTioWnZwgbgy4ve
nNW2y4YdUh9MqG4Z2D6uQz13wzc0kvTP0CVkiiQ1fZEPS/sk8YM/8WveTullp0wo
S6yYT4j6yObMTfKnCFXXY4Zgdp8uIDi7svPxfkDmybPhFxoK/L+MqShIs+mzQ95P
V4r74sHnqnFrOZJ+D5nE8RfQUsaFxlt/IWgU15p1mWMCBR4PGGBDvbNYbL6+MX6q
aAJxQHFbqiQYNnjvW2hczV0K4lm0uHyEyq8DQmUpsCu0IjEHqYovv5bEi0L9K6eK
L+SeAAyWlWq4QO4RGAgVQ99buPEhoidbQR4RKBIMMcHA010Ch/gA5LSGIW+/8XK3
xY/QDzfvuzmhDhIbKA9/qGAUfPSUanIdfCf9aXQ+6TQXJ2NsAlT4TwzSItu7Y2EG
F4+jKAxeTIHc2cOURgYR7VLWZgQqOEIt8ZxmSLFZocrltC08LJq4AkZ+WF5VkiCG
pqi54nGUcvZn1NoE/YDLg2MtWif3AqseTyKM4g/J3dzaJ3vUrGLKuwwII0nDsIRw
CgzpstdEh4xGE6K9fTJhgsLiWZ443KzZR2+A/w71CSFWqZQaNLznPOfYBKTOkxKW
AfYGmZwlHxfoHgSypaiptdPBOgDYHWmmlInAod21abQO9C1ZrtC2FJ3LKZmjSayj
GJVfBoyjZFASWeKytRGEQ99Gbu5Vh6t3OPWxv09+w9NV3VV+WnFEo+ovbqUO2y5G
jkc+NJBHAQQ16BhbciOp2oayus2oD2bO3lQPdaBHLoImXVxe/nGqojZ24KtuLxTj
pRkC5kyuVfXy77xr3Qnybo0B7PuKnJv5Z91g/4R0oWs5qbje+pcSHLFJYqB1shMU
R48Am38zP6usL7gfv0TlVe3I0KYHmWV/WQyAWw65EVVZaOJtT5Er9DUwvPwitLib
nIlYvR98rBtcENMCaY7B/qxczDRIlqoN1lgBKvhRKk9bqeu3eSl7evzR4Y9G4G3G
+5VXJ89sfIAKClSM37uJ4zDHhPznDlMOQxrtGKKjbWR3NwopqU5PvYULmn1MP+d3
LPUXVqfg4jECsM3WI9+5ovurfUN5kBteUNC27k+V785hrRIWHYjzUjD+4a7Czwr/
WwquEdAomdls51Kal8kYASvQEOEXm9TCRJGJyGB3isxvHS3Yh/tFydeU1ZCbZN49
gWdjtfzKGzQpC2/X/4wBOK1FnBr6ACRAzncEHFBprbJAxk0R183q7/HgZhM6gBHW
B8ipG398ngjH9Nior8/A3jkWPk9EaANEWPPYOyAW44lZIK24R5GOM5qXCWMePrOn
yv/kMOi1povLRkj6ttrY9xXyojh4VZh39JGvt2ESEf9U8zz+dn6uXbQPJ5N6JVdF
pXPgXWVDi/YbM1olUimBKSVItxAGXLTtnWDimRZMwcSgp7c8qP6BBce8ucnmCtH5
RDK0C2hlfYrPI71h6WHb67j5WGxuDxOnYBgWabPCTwlKVS32OJM3iBVWzXkF+Hv9
JJqaJX8Cy9sqCiDh9L2O+8ISCw29PCCGgP6P571Fq8SIZH01TRHzKayAOGCidrNc
mU9cMpHE+rr2DefwekRdSH4YEd0TqvXxV0xArgWOboQ5zdUNxRVzbg6IWpIfIA46
pzlhid2qJm9gINMIOrYmlOaOcbxobTEbq+CyIP8rgXzTpjXhVckCpUXRzJz2/vRW
FwUtq/19CGMNds8FR+JjaxXJs96hAn7D6valq5mrKDxOxysoguQYIlHJ138NI2vj
D8NixgVpQ22yZ/XAkmxRImzO76AqGWGa5ARLxFLPGNwfvS34KJuJK94aBODXSGoh
ghqqU+b79A8TAR9apH7DZZACHbnWx5dlhclSDkRLUbJEKw/D0O7IAC2fmC6h2Pw0
gTbI6CqXw46F8akASRQlSs92JeKgu5dH/1X3VLJwij8cKxwMGyGxBZPqw/DzV+KL
XWOF42pZkIb9KKcYR2neaiAcOu0oJn4W1d93zSs9Y4bnwu32a7LE0qJWWV5FiCLq
JLnHjM8ADjnkPmxPyADF8LWgO+dYV9ZPzFDMq7UDxKTYcoqc80qU5ODu/fksyF9F
bzQ2wArq29MSgQK3Z7pexvaKFWJk1w7+unUAJ3Bu3ci8GqLa5tVh/ll0Hs/l/+Q2
xHh+ncgIgOjj4i1REKKfAp++gy0vkKPuw2j/ro5PUZnhuF5R16Eq3FywGyNPexpP
Nq20cBjgN57sH9foH8gdHZl10S+m38c3u3tdy046bS8lQfadVwfrPDJQKF+scY/O
`pragma protect end_protected
