// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LIz+ylhgCU+k0z+lc1gJbJKCdf4ss/hxwkqiyUh8leySWXGp2rgwtVupRpKG9C83
gYwszxE31LUwhYnflgLFJWbfUBMA1OMsS1E6e1yUUJemO9bx8QUeQ4GP8MAMQlcC
7qbp1/AfPEHkcOhfePptMSWNq5lvC6J94mqeRa8BmAI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5440)
u832YUxMhQKR6SWUZKde84h1oXrIGcIbyvheazTi8xAney1uA3q51vsfJIZyXZaQ
DPCrWcAwojM9raftOnXiODuP3cbvrIwM5gxK/N8kv32/SP3yQgDYznPGorfMarP7
artKBJfva0tpynvv0Kclg9WZ1kCKuL9DmbGQtNLE/9+uxkDi0mc1v/b7oyUS78s9
ofpo+UQTJdnCgmMnWnCbwV2WVG6jCCkaYCM0/DPgTU+MHsdJVCT9fsLIZgzyuRj3
aKlkx2CyAajkHjwjMg6NtFkNgEt/3Bk8RjPZW3PNoFA4iZ0oRot8Y0PYk3d4xDlf
QLd/xkTx5XNbTm/bemoyvyZMkwFTamtVrMUtpgdYAQJ0ixkzC0ISD9qQbfYYU+BN
GHtkbJ+4PgFHzrxoL4AqK6oUx46IfjXmXYnB2/Jtbymu1LAI33ivaRolKoWhd5aV
Lt4ehc5UWyACAtYiIxd2ErYSHFZPgLK+ocCqsur+1dSdjpCTxIfjtbjYqk/gvZ4C
hr4QbrhUp8aWs0Gs+HliOrWg1emP8896RifdhEpdOv5nMLeahSC72UxW3JDxeAy4
EBgE1eFF8kSsQJ3QefVZ4ZmO1kyj5QriaryMYMBD0BQB6LubDdLcrvabKOOBiGIc
VCMpOCxgREL6Wq92G1kPWiokTNpAc8p8ae6IIxwiWepG4075ePGzqzOM+sNo9TgO
TZ9AaJT2Jkf5VjJ5ybyO5NmHq2IzXCIuINea4YmhwTdSN91leGobLf64wfCzxl9a
huEFCE6rjDb3BEIJqEw9+Y+Qa/SBzMfDL/Qf9zzYewI3ZkBEBGjTR1SU7td4D63M
clcFJxXwKMDlmJD8RQx3Tpiaq/cxdjQID3P3QdpDaTzTmS9VcbYt/NIuLDCNnVJn
xC0P+Aw1zL6IoF0/qhoBPVTH3DNC2GXz5zQZSdeInkirwoyx1mp+fsf+K89LnNBu
tdnMpKSTs6Q/XRmvNi1yetzA5J07dT6f3faDmr8z99Caf6erj4qJQLkYxuQMNxyo
vOTtJESz8D4T3g5TXCE7ALODUN1HJSRcfHouveXEswzcgIZqSwPImdS5j6hKhnVT
G0/rXZA5w/VNJBnyVkS5dKwdRjXAcmlmF2VeDIb7hd/A61BWcLULmi5lscKNOY39
eDiKKsiQJ2J02Uk8dY01APfePAPJbhfZQQG64IcRPzrJ1BBlKrsbUwKayOIfdFPl
MxuafGKWM2C7GQAz9QL5rYX6jsCP46bnwzUV1QzL308s3M33qFwuf61R8VC979bB
DCiLcWZO93SK6gICyDQVLZ66SRCxXqmgHonK3q4qXqizOEuHHqoueCFvcPS9CY9p
b/eHekLziEYMLBFY70+MQUAUHV4K3U/7hOCMjvGiVZJPXeuYvN0AkGBSc35t0WEO
Hud459Hxv/mR9CsKiIJacchw+tsq/FW0xl2ylsgeUt0nw+qszWYdrg9LmGHcVVrr
kgZD7q2kSQhlY2JPDsIDKmm27RLiUpMtnRxTFdDbWsAQNRFoAURUIBFUAB0wDbKl
oTWVEoEGHS3ceKltTvRy/SlbaY5wZSM0rFOXPYRd0/atO4+awYOpNAEXayM7SZ5S
xcoFPF2ISpuHCLXNV2yY3feCWeAd6Wl+NcXbzfGAN+B5mjslhXEYbhGR7E5PPeLl
1sa1T+JcWnpqjDnmVF7JlIieS5YorckVhjh92SUuwQ8J5u3hDOhbIFpSpyH0/Awy
GxsB5ouCcp74Kep/dqeEsnmd2DNoAzeO4mTW6KUN/r8TfOm06D1UTcmE7IyenKEI
h8mXJaiAg2FX6WiG41qjEjq+WCBIxLzhhaKbp+fh8zFDvziq/uW2RyMyodIstL56
Y9p8O3vPllXBPwJ3nQEXSPWubLc8rIcEqotlJeYuIQSjtnHuhQ3K5iiBc5HSEKB7
/ABjFRRkOxOnw+/vQGdbv1A3yisYtjLuwMRXsXrNYZXiv//v7mEogxWSuEkYYjXG
igds65LnfMDrN99BJDXFOLS9B0mNQAqX0jqZkGhgq0SF7pCq8UedTf65DM3iTMdc
8saCHS7PQr/9QG+Pd/lCBnzAUZPfy78YUCdkZMQaaeYHFFKts31GB+KP9eho+I3X
8udW0PDeUZ+WWTE+9oOerNkCpQkoS+80XP6VOpHD4l+7wiOxDEmu+dc/QamR3HPQ
TmRj/CIG87N9cp9wVjqvPeXUWgLsaCov4EJSBf8MfxEc4fe7jDqkJEyHK/6ziudn
SFBowf7JD4P4Z8YEb/2Ukz9RaiZEIeqKbJ478iglzrtRNq0+N4NVzmPow8y4cGYw
c9VXsApBSl4YBangSZldt0NJQ9EjK8F+bObAjibyMn8XBI02ZkDgUKxK/1plq2NR
lgmpXpuuC8KSgkcH79FRnXfkfyp25lMoyFRD/7Xfn64TEs14EJBolbxIMOs0yh0Z
I3/kg3JYuL6eaEiT4VESHFZ745Z2lVRxcJ4R+uNWPGTn0TZn+fDJ67fusVg1ntiF
eAfaYF7ev9E3hsPzzsqMwz2xrGhi+Nrn1z3DcegbpOR46j/1aHOYyxmsLzm8rPez
fUb9ZIVBATVDRIjLdD+kGB8b1dYHWQFt/N5RO9/e/kwYguodqGxF0siLMEuLKSB3
9KWd2HBx7fchyUtdKOxG8bOZWxvOvVjnS4nvr26+KV1sko35QRruH0F8rUs2Uu4Z
9xmhgLflOuCXcy01ERwDTraP4I0/zyZdtfTXRwRHgZW7lnGpwQ2efcPZIVuE9A5p
gvfsjNJ7lohNujILfSXCvrJnwK9GDumI1e8U5OAcLUNl96yKXVwuWv/NqVLaacNs
yMWu3SPLa7ZiL2WK8/TPg3PgJBjCu+4sQVRYOUBsZ7NreMzqXzp/DJkMWLwfk6Lk
S0ImF0aEqR4+MDSxIpmh++xrX/G5Ylx+dgkWsp4JuKFflj827e7uUcyGuQOvq103
IBG5FvE3AtYWDuohvL0vnkmuotGPvNSmS97MNURAAupJzHuDhSKCgKvs0/eP8B79
/aABCdNfdiePExl1lBhGJoXkmja4Xb6Lb7RE1OOoRure+m2ctwLA2fzoECkyyI4d
f1WQVXYp6y4HyxxaQijyJ5ZJuSNbm0RbhT31s5Ytg1Qed7sO/+kS9Iv2xgCDp7aw
A5N01Z1NJ8Euc3dhhOCFNjg1Bkju6Q+NJTCc+B+U/ITO7IwKBBb4HBhenwTECEWv
DH16u/tWsbGIsYQJLMQ6K8+Fv4dO7z9a+q/UNk5HN9VMY6BOoENmQWNIESwj3cIk
fop/qf2cd2AfE+B6UsFY7FcjMvgdKlzAwmoFE9Nxvn+qRqpj0Dd5vlT6HwYbcdF3
CFjwJAJkI6IgaoNRr70cRn6BiVNkN3n5+B+uQeubkejxHiATA2mD6/fvDQj5xF1u
4al3MUnvLT7gX47Y5XBNYcOsNNoIXha7z/ZSTLd9kOqFeY2c4DNSRZJFENRZkR8k
GJXByli0yjGZkbRyG2fLm0tvISabTSfQxZVx/hjrd4ztM8Bw5tLW5y9aJ0N0H1QO
OPPDhuQiFe4LZvwxqwv/xDLNjYd3OSpIGaFdFKhfaoIQZ7SrkTTzCQl2fFzvF5Qd
wiYIP3tCDiZ32HEXAQm57242cTaJsB85+WgiD3wGmXVfXzvap3zroqgjohWQ2hCg
Q6wqdCRcY+M5P7aeQFDItomS7jjaw8Ev2FMMEMWySYj8sXsl+T3gC4neJkSNuXpe
XZ2zBkKseTMk2rRiDVZUvUiDzPtVo6hqj2t3vXtLS986OFU7nsk6kRcvS1gl0ico
3XE7yjfsAQseOm2/s6pqwXIJxr3ty2AwqN4KuXUS0SJ79Zdb4PrT4a3NeIhgtil1
3AD2Bv6xGT5DzbzPWgc1p3sip4FZ5MaErRN9oH1YhYUC5Uu4CvXWGs3Hw3NdaxT+
IQR0Mxop7cHcxI4eE2pNtZU9IOlhhvKAmqDMfsQjJZoXXs4kt5T0K+denhXfUsFJ
j0mL4BBpnmcdc87cp6Tbz/6y3Y3EUiwIbuSz4p4pVmSMLps/CgIsPXsLGpp+Rib7
lSgLh+92otR96H2RzLS44D+t6YHQkSFSm6zCuzjUMMLJlkUmkJtd6OTaRJgy34ex
wnp4ys8ppfJ+jAVDM5hV7tzqpy6GMReJrMkDDIK14WN0aArq1Hei385HdRerzeYC
77ZO2oEDfupoO27i4cdwGwGBhoEgxI/dru1Fg+qstt3g70KjrGRGEthgp17i24UK
Y5RV1Nk278+ZkNgv/R471ydo12qz6/Fu9eaapD0QDxEoKzcG8ulVvdwI8mRMVv1q
GHmRFfgGlhE2CReKo3iZfET8XegJnZXEY/0A90Or7+V/e4umRZ/QubWWtUsY+uj8
pJh4itIboj5TV0Hy4FKfF3VyjATfaHKfjVfr0rleSA2PZnwkaMsU1++gnRzNLSnB
4+PCug8bYIj1VqLbaaBmfDBvZeqGYb6Jejub+CW52SV8pKy0rvNlZhMOpOo+a+lv
oxEIZ6We9erUW16lw0k73HbZARNcdMHraq7KJjDEmln5mkebEQ9gQD7H2SL0i3Sw
zk14ICcelEesJhqnAD0pz97x9tu8orPNLSDKhXmHP5Wusfyf5bCD2yBCAW+rTGUb
zUZUmKwx8KMeVYWGFo5XOqB8RLymbx/+kCkI3joUJ0bcw6DGKo2oLLnnOhQHVM3Y
futaXXKwQQt4nTlPCbqi2XBG56ZTpZAEuoislWe0o937pYpZ8wL6ScRMcI7T3Wog
++BezCsTqcj+zUKTECeobX0S4DVYa26ucr5zyyqpOARTzZmDtrwX/CQFBf4NN0nV
3vwNoHiOWwnsBlHm/q0MQLZ51vXAXcG2I5eXI82350pKuKjZXSHOQ+ILPO/4dk1I
5a8MJXmRxHQp/hEocME1p3oyPYlzjvexawmMC9jGAGcEWEgKUiuEzHymaSSAAaRu
XlPysxNX+x4m2RrTlCrTrM/6OfyicJUrPeJlHXgoqecowZY0oMr6Dja4FvDBVHFp
74mtEfHEjdboBeotU8riqwvcG+Kn9Fqj2pYuCJ22r/c7gz0Pa8jVeZ/aHFhiekUI
0R14bfAQbg696fIK6ZSfaAxRpLEZ13G4GT0BtessuSOKRPIrLfycPJuG8xlemDxJ
hVMvNQoXbl9FP3GS8GFtzLtUJkUks3gkTINTd0sx+T8HyQBSvLoBEu565TCItwuW
oeQNeuOZ8nBMquSzZ1h/Ui/xvMtUHySbTFqEaDgslBH/JPvEV6fi6BwzkigVTHwP
Sf088FHjUOb3hQU3vmzm1WnICzFaqAC1Iq+4ozfnqqR8NTvtQpmm34c/Ku0GalNz
jP604VR6hAXe6JHGD7Gbq2naHfGC4IRwLhHdGdxawVD4Jid0EenVR2CBNcDyZKTA
+Wo44OxPWGv+Ho8hp0P1rY/3Nsh6pzf2feln4dm2h0mJ6AYiNirC1z0b5PO9/sjV
7d5W/5I9zRTRsgsM4DikshpvnSJyMsZc94zLvuso9hICUA/0Ped7AFRqiANJvcPI
xb3qkuN87WJT0lrhtCihgZEse9cKxf1uABFsGeaEBM4HQlqRH5ISAlstcS15TZk3
nTXab9VB106tyu1YYNgjvUEz5nKXbFt2YBne1sqSbULG7/+x5lO7xG1yPyz12PFY
9Bhyl90EI2QyRgBFe5hUdLpEfblUeZqnkodQgj6t9y70oyKGUr1LsaLKxem7xOOj
XxMvpbWATP5Kb5A4PWT6NNTIkccQhkI5ffx5XhDCZWmRw8r8nTXzetBmRHea66ut
PtS7HVpk/A3LEeC/pB2t3W7S/24Bsscs4J5X6QNVSmc6R97dMjSMADl1MAAkDytF
6Dcon+EcxeveKuI0s9q1pKqpogSj493c8Tdx8Pr0oaNdTQbbsavWIj96ppoAvjsZ
pPnn77p7lwhzU278x4lK6MdY9d0cjj9VgWbpQKev/Su7ZGkiS12ChflkQLUOb7Po
aX2M928wwnLQUi2Du+SpF42coGrFhs2yEbtsXBIzEhbXxgOKRRSJ+rU62/qIigRp
x2AUEFl/uF4qMao6dY4eEEm6R9tIUkqijmZNQOIqsLCkNah4XXik83HNBpp/nFze
PCGfXUDqrPuQjtKH8elMNA5Wz3XEYSDjqhaF+0/JU+dzA7cJS5jeuRP6XjD7Rs/U
AI5f8e/XSSkK4OZB9qS5wQjav4govcCNdrVeTaMNbR6H0cxRXfHXFsDzgJQsEXou
qqt1+Ajz702sQNVcDoxpDOE1aLcsnvt6lCOsCTX2LJF8xlxdTCyiS45ekCmiUWYL
T7QJ2WIvV0QaoEgNk6iarLg82kixhM5gvStlA2biBfQb9l9MYgDyDbSvHB0vs5pw
HuXRur1uB1lxuy8I1rD3ImhjG1qBLj9GBOwvf0LLpAss9WuGnzj86u2jdS/cVqVS
Qq7pERFajz+r6oO23xUFdDnoghHhqjIkcusF8KwtXz5Ak+oV7jO+UNrNIHq7aQXm
3Re0mq2+AdYEr4gBGoSmgN8I5ICmJqC2vUapQEorME2+QaC0tU410xCBCOnuOmF/
a57vy8+oxr1Y1iEnjv7uqSlnqa3WQhb4lQZnA4JrwL/pyviRS6M/q3nF/l22uLzp
7iTyXcaxADzMgWPmaQe0Q5Yv4Rxpm1rHpKpqd8J2Wa/V3fWDLI704dYVc70GGRnA
c0j8kC+AOBM86kM8lbIj82mGImKHg2/m3RSNKcaCPcETFzPDKUe0pfHmMsoEXVkc
OqjOR+mJ6WP6/paeIzEpCQGa58ENhZZJXH5+3nBLmrsBATZVtYQHqF1/QdYIP7Uv
6qrXEvVZZKEfLc9NFkGf5UrskmxhiE2WmvcwGF9Rk6j5q8yJSHD0gV7BLC7/eqBm
6ecWnzeHjRldziZLUhAijEOOA5SCfa0FV1Hr14ac69vCht08YVX70XhLtaLYsItm
olE8TVsAMyxEWV7UA4rc2QxofBpDqQ803iJTm7J/PzdL/VGoD2EU05HEhrcXjwxi
jbsGDSBf/g2Q0aaKHJaboVXkjuFtmL0hPwWmpGLEKTMjjkc/uujkWatTAhec/2vm
n/IrjMUe4Upb2rI01igs2/V5zLL/cTsEoeEo5o4qxBiirbb4uL1/DJpQPdWeRvdd
KyViZaeGDypjCvDlDKjX1jnksdV6hadQouRSy5PysP+RGvhX1ajslEbxDRNr4kAM
r7nygz1OVRfPwShECwJ8j9QQSyYejoGuSzsVUR/tnCxT1sCm7HZZj7ML/Uph0Nok
mcm/mzUyWAmlejAKCC8Mxw==
`pragma protect end_protected
