// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:49 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E7MXIHV8WFDIJ8aXSs6UZ8ERP3I+8XkDqcP8uo2/kyAtOYKazcLhTVhkT+z8RvIP
Np5XJJdEdj3YhkJbwHGBjlkF3+Tq7CFJGbvmsv8WpPbR0YryG/0lKMZ4PDyAgUyl
x49DgaKN8LCrXX0CMJSfesCrWfRhpaddqkfTMXwvaZk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2720)
C/U9kHO1ug3V0ywOrTEsAH/qyoJzCaBzDrhGTRakoUzlLw0MutnHR+zBw4CDZZ2y
ZrPfs+tQa3vyfW9qHkAhb4wrly7ez75b7xO3GuE/V7gnRYLol0PORCYlw2JvLRJj
TTE0trqvCqvYPqCSmO1eRWhqYcdXGTcUssK7wzb2j87p05tJyo2Xvz8L8l4HxBns
EnuMK+jd5IyGoHHfnruLzVkGuTJdn5gy47lEpk2ZFDGhXxtLnjAOdsNN6G4u1Qii
lKq8AwKWKv1JV2fTGy+slyltlVgSpIldLG4fwWdbP1RM3kVk1q+bkdZOh7yH1PsG
bS4wOTDMLLW4sQYnzvU2VMZ6U1ZMA95lGg98Zj83qMz5ymqeoiIvlG8017X6Kxyl
JjDcEHMrs+z0WBinB2eZ5AKDD6B8IaGgbxEipTNLnONZt4IkMoQ9WGIQyqDL5quB
Lfuy4DPOFLFINit/EH41B0I0rXORddaMZaeUpyp56JQoND5JtlprpyR8SVlrc8lv
7fLm6BFjI9tAmLMUudghUaG77pECUFE5zlw+WZ4Luw+c7Vlp2G3/U72NDsxvp3QA
r+84clQuEA74Ck7btaZNuv1FiCGyS43AgMpE7NkA3nitSKaydJ4gtkopLq56e7pq
uC4LjkebH/+ir3PuFSL7wXP8124P0zxqzcZ8ZE9RB3R2eAla+2xCMeua54Wi8d+6
fGJ+DUBXcACn0aMcsE8QExTInX8VkHA6MMqJMzrsZvq717bH4aWLnIlJUBieYpe7
ZKkAxLxOYqj09wj2Dvcbukfz9tj937mOELmX0hbR4UEp4OREEhYiSrCeEKmp3nmA
eazUoimwe9c0ekaKtvmE2sIjpRxLomvAzIdQtWyPy+HPW1HR/juxMvbtdOcfHji0
+9S8XsZQEHGj5oC259eKKSvl8ej/b6OA5oYtR+8vDm4W7jcr1eQEv3haOUr9Y+dS
GPswuxXR41emZb+L2wsfDLezsNQlU3agbLjSERsowGmo0xLSIEb4jbh2rlJYMNPP
rMqTpJmh2IjCGBpmUMBUatRY4T6K2P38LA0NbjXQ/bIq3agn+kqpiEPrN5DTq1Sg
yG7R1vTZoind35Ss+mp9WrogUFxKwPu1q998GWfqjAgNUmmQPgiOy6q7g3CUQk9L
A3kfIULlKQXqdzXCR+whnPB3hQKL0zqH6JckO+TFWSiphihQEvLMH5Gt1Ukeas9e
ELqTJiSla3krwvg3MXSeofIibrZYSvqs5fRZ3w0+hnsfJ+jg3EiP/NMCbRtiEh/O
U6pj0zHN5QDzXSTDoVOiOVPmsUcALSCVM92cEJNwAbBp+//Iq92Vywbnzyv2jvg2
aJhtmO/Sw5XsIDa76XG6uE2atEXTqxPdpR0o6YfBX1yLgX2DmwZByzF1RUT0h1ER
VkeK6PxGMKWX+KU7GJbXberRpVFIeUQo2C+ZshPC8CVwApqQzDfS4Q9Bt5+q2Fnt
8R0ij1CNSdIYxUF9wqVIBCaWYygYd7deiV7ggBVdO3d9gAO8GCenemUP31bWUHvT
QmOK08De95hK/Ie3q+kgEAZIwY4R8j9kMk74URQeeLAeLXemdUZw9AwheyU/uq1X
dFbU3yF+bf1zUuvOJbb6z9t+2HEiH20WIoGn3oGChlFEUyd1FkoKtvIlzTPbzm6Q
Oi1aZynvC8c5BtJc98A2kxqZiJb4w+8lKtMH56gIxSnUotI//o3M8XLDcdAFoHD7
f/le5RBZYwm0c550tTvz5k2bqZKXVbwhcisO//b36Vsuu7tQjPfXPXHsqzGGjEsL
gGTfUk8kQLUcIvczESmS/n3kk0YTGF9gMqwCymUdMLu+xcGJOPbOAfavu4uqYwMB
kXEYzv8xNGeNrmnz3EFIvah72dGzmgyo5ao+WOfJ2yhMoaHROOGSmg1TmbcpIlBX
ybestXdU2Y/bOBlRsGCjfarvgJsuv7W9ISbOvdelZ+zLkT6ejBXtzvEPJu3izN3H
9pONiyu0IDUmSQcgrOrgBNjL7VawtArxCRiVNBcMW8BKEX80GyGdUS4Fa5gpMPG+
Re6eKEElBCnG3MYcwYPMhUxs9GjEFMEZaFBFtlCyOhBWNHg4xrDW7v/AAsI4/7gg
+QyX94MZY9SwUlC6kCAsgJzBWUL1Il8ikaQfRgjcOckH2PUYTZ4Z2xYzT9eXXpb/
ybeyW6fazYg2ERYiTNyxy4AbyebX59VuKfyIq88H/ClrxiAYcrPxCq9Oxl5AWfIh
NnNpy7m8IIFCvOlwPG7EbDkbjffq97zDu3CGa/Jk3b+rteRvNQ0NcRiZD2Ii6pC/
Kts5GdeVU5x1cYLU7KqKgCEHtGWDBAUQ1cc362xSsisyw/mTn71MEFeZ8WiZxD+w
ETO7txKsrC6pAFErBftEy/0gSWG2t7DbXyI6ytWcnDmyzv9GdqWi8rWk6zRnaGpT
yuYHFyyJUYZbtdRC23CeJU12vF/nH1lGGp2SlRTUbFfmMz0nb/nkYJIZHzEgXvOI
ZZjF7ibkTfmTedfRDHqhWAjePWbNRpjM36A98+tKEwE5dTyBkORqb5tgqA1NSdrX
8GZtyYOZLXKXL2bUR7iEMNi2GfcfAC1Smvdr6GsOLoZhPvk+UHTc43cNTuMlzk//
7x9lykj+EYSvso1E12p9fBUmsmNAscfH3CQMTkSFxaFy0wDTBBTTA+n7LSmj87jC
U1ODDE64rtxWeG0NBOJ1u3aexNkNaNJRVhSUZvbuPxQNJzGkQMCQiy90tiifOamu
7m7D6eLqYZQdBsF8wVaQfEX2oSVFFarPdOQDb3/4Ft0o2T8KjfLC9fnynZegF6O8
GEKzAkTHd0APAC9+X4cSqQzF9KxRx+5EPbM+QvPgobbMYr2/K310a6ABrPspl52X
J08gEm0R/1v/T0J4beiAbRKe+/x9DfbXZt/iYLnHN6U0jI0Swt5gKdyrCzl8GsPR
uV0FpolV4bMd3KtdJC1eOGsMU98EfsD7o+ILEgfXqIYxkNSS5aNDhCFTU9aaI55l
hT8KNqhBdBiPrOnvNACc642j2PXxfBwRFkBsuGzxoJyA8sgQBVTUG9IX4ng3MD3V
MknJjhvhhszBJWdJSomVxtnNeAeEHZEAJIsuiQ23RfnlmLhrukzn9hJlqn7c1qzd
Na5055buaY3hlkdY9LBssmc5ZJxxw6by2qI3O9H/nfSAPnGkXiVwLw7a4YepdXDT
hFBuMeJwm5vPn9tsNBwtEy+VIpKImt2gcCZ8WPYjOhDZKKX6mhg2fcWUH0yB0WMx
HvHHBTf7KZbeP7mTp8S0ChffOuQUsPxct5YF91CroozaX5CAlHXpBw4i+HutV9E/
jcU3QWAOCQ4hMo4R/KHNzALjtZ04nxYnhmGbEd8gg7d3g9zkLS9uB7ETHKISWCaM
Z1JdYzo86c7YBc7EbYhx3+qFBR0FQ9RcfqMF7G/TgsXnlfYkPETzUCuvfG9dUALj
O/xaYgayYd9o27xQh736a0lh0i2JltBwNl88jTt3PEilMFqp2JIBrmVLxl2gxdS1
M1QN2lIjDfI35/Tdwg2AyMqXge0XFR29GY9boFnDy7eSotbSW4Fcavx45icP+ObZ
TJ45UfDDLIlyavwhMd86uRTOpFjH0vhUy8PoXj1rCUY=
`pragma protect end_protected
