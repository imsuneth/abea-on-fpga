// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:45 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Snodm2YsljpNAPnnt0EIduMtZjcKAX8iKoFteA1eG6+0lf9HoPGMHU4k7xnj0qLV
H70jfHyiIfMKuDBeMZsOFJrKXRKbODqp8fIJ7RyHSaW9e/dIQGQbQd8pDJb96667
QxYGZbiGcD8GHGuEriuQ6WyThxQTGx0HFMWdLxpJl8I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4192)
jAwITbgU0HZlHXZW/rQJwMJn38sBeHhoAqNhR4HzA5PfljPvf4PQ1NzYVH/qleve
dcxqOA9sZ491znr1IhjxiNoJ21ktXzMA+kk6202WZSwM38OIzoyD6VrXBQIOqMKG
oxn1XkLfpbqHeOds59CyLqMeM6VX7ejDnzqmB8f0L2Y97snxPNFVTmVuGy51euD9
DKIQJNj7GU4ofwywZ2vjFNmeq1y/4vxfdzXYzWnjb2LU4WN7aye3N31g3V8+noLo
2O716RInX7uLG7FRB8NmyJvFPYr4AhqI+Oo8MAyVa0JiK0At1vokSPvmq4e6W4C2
VGKUlDZghqTXJpYacm53SYkAg/ZqiDQzUvAbjbPgDrNqKCLxFZrLKf9tEtPns/R3
UP1KOwf+zVn8ryejP3inTcgsyElQNKPdlzzHbok0I0eBwRvnW5uiGnSTdZ25dmMc
ESIS7Y7z/5pgpQBcZ56iDcCH0Mg6HgK4PGQP7KFHqagbUwV4ed6gBDv3PiUUJdzc
zPPgG1fl0epi5LPr3vp2q4Pe/UKrezILPvdX2XA8i9t4wivW0dodNfSQgl0yAXVZ
/FyeOgau1nnlO9qzfXSO/W+ThlrxxFGhUaFEVDQazMLaIKXRWTWo/2sG3Uv2WubE
QYdA+4Q99Wp0NcNPmTn/JFDhjj+3JUD4ByfoTbhrY/o4s3g2XRa0CnD7JzVfhjg7
F5ZP9jSPOXLG8av6aO6ubLszqXf1vVG7dvV12BVOZ3XCycJzvw+MXx1Oytzdppb1
oIVz46KZXaKLE6XV8ipfKY3OjM+d2W8/iISXdvTrqSY2uA1OGkOGvPG5SAMt0mUd
5Zm85KgM5xl49KanihB9IcPyYAh28DDOvYSWfP7YcchuFDASWK89wm8qwOz71l7/
VVCDAvq7gywUD6nzAcV7j8gIKY9B7Kj+1pS3SR1+DV0rz+8Xusfr494dEZtREQ+3
pn2fVVg0aDyA5008Eo32Qt8WAf7XzBMOmIWXzAYSsgfsIn6GsLxAiCZwJxxhIrrC
Pb4ePxXXyZCTXBnae8Euy38ekKod7Opk2H9B7fM0BMEJbWTCZI2GgN+BMZ8UyWsB
NycNIIpD4WTnbibv9Xin8v3PLtfr5tNIO+TDb9jRchrR6ygNItXjERJYKc6WZp9x
MG7MetMgfQAr8iEbqMfLir692rBSButfFQPr4LvBkHhv8yC3mfVMExqyHNLcRAxX
JW25WR3gdJy9thB7I3XsTRc6efn3yop3O6ean5LS2yPRZOo61km1hH7QdiSIxz4x
vlvHgrTCC7f9DWxZzbWIAiAkBpBnSCsnh9qe+K099pgbM8vgYc3377K/KNQy+jB0
QruKf+cIog6x+cA/1MX5sNJGaTKlH6NNqxzWo4bNBtKWwLOwlmhPB7WcMpfxgsb1
V2qVdeaYvePQ+OPYLJFzyiedB+PbEhutVCSXB9b6l7p4Jds7hqZKgL+knS51j/pc
k31L5rCbAOOh/xQjLUgXtwNXPJ4xXSzfGc6tyUtelx8vds6+eDVCTvuNYN3dPya+
g3xqiOz98P4zQrCxjMxhptPj9zdD5GT1uXy0lHJ3JjES40e+DHkOVkun4bLvuoSw
oaa6dsCuvJESji/I3n/2fMlF5XjOc973Ba8PlvtYWk9lmpRaZhL9CRl6tIoJ34U9
hPTmyeAbugpv3X4j6TE1ShNC0c0U4G9E5PohaQV4dGyGweg1sFPQiKCdH+QEH9c/
LjYm+lxJWp+ks2X17kAWPy1h3b2SbLBSORfta8yWjcp5CEASSBnBGmAWlyPmWjKe
zRsVC9wXtHYP/mio37cENYF9TzTlUdh8q0ZsCU071bo1hnNECSxM9vecWejXy6HF
5XJwgD8Vu2FzQWHOXUFwQ9uM+irbRaFVjym5Dty/IP8s6cLdY5VxUyfe0f/AOkP5
f0MYQ8AR5VwKTD93xK/EFvbRs9/j3LA2UR3u6JtDjKmDnJRjsB8TgQujMruPjhw2
tU5r3lOTkzsQ9wam4NVSQigqvjGfGDhXyY8kWCBv5WeMmuqLcfQ4feNwjOeNCWaJ
CpoW+RUMzIqB7rXDHY2gRwzvLBkvTf9ekpbdqidAZeXFnB7mzwJasZGam+9ZABuQ
Yx6uFb8/aUduQyJ33BqqeyfNwvSXedj4eBf6+BzONgvlEAEgvEvsj9qU496FEGh1
BRj/vx4a6Ob4nkm7bDQ1csP+ydVgjx45UZyF0VvO3ykbv7KdkBs82gaJapcZO5fQ
aXyffD4iuyPg9lHTAfcbXGEJYNvgklt4wAK/j9NfbLsCZcWUcuKMcOVlC0FSxxFZ
T1WlCx2r7eja0yf+sUPZcpPhE5xLDy2thxgxF5fTkUhybSYLJFBXGnRK+0CAS9bZ
Pl7G78DSPILjTYKQWxwv4wRfA7IYhho4zpvbfG5E2uUMvAXbEsZ65dOUy+IkcpUp
eKaznZIlNCY/dz9OkoTOIsPdV2XFMizoyxS6htrOf8LxTpmBaw7ocJs/ghvh480q
ppD4fTIEexkskwPI4QJwPHtqvQsqft6t9u+3EY6TMeJ31e+Esr6nd23jn8+kKhZH
OdGRkggiWPfKbIrPxkTpBVs4KeOxtutLEfyEWUi3REdGLADDGPnk01I0zACOjmOb
fG6Kdz27EG5bMXMoXrXk+J74uodUuE96dqyrM4lHSNNzZKZGGcvSgyfL+Su5a/5m
Qco85S9KkuEXk4eeQPX1HsGNbdveNOD/4OL1j5c/UzG8cPfnUdgXXoDIJoCmhGbR
5oXDr+Ob9JmfEkY1Oh6I5Mo3HU3MSBITNenOJkTAoqSiOBZkrBLUNOY3AEWy7AYd
HfrsaME+ln4JJ8eFsKZwjPs3lXiviH104zojKkd7GzIwrMh0R2HY/McZ96pagjwU
rA1YRE9waSTp6TSn9gn0Wx2xqzMtKDtotGLvEy5zlFGORgA3tbM6Mmo1cn8Nkg0U
FpncR449nVgTLb5WWRLia9A88UJkqSWWy8nfMBexljFqXNb2Mg8GkVm556cfHBgV
dIBEx4EnAejOJPZaY257U2k31Lb8N/XsFzUg4Nnf83d9r5dtCR+iTUvxNqoBb13x
DEzeqFOkfeZrqfsdbNrt0VSrFNMcusACdVvqgYovaAVFAMKxTB4+isEXliTIFN0w
UKY/Fj2ZYhi+GjDKBW/anHBOFF4hjnNXViiD2iJid5GgobZGjPZX4D7gfbdY/dhd
mgc0Ta7f4WmqQs/pKmVZK4GuAc7Pj3Vz1Lc6gQ9Xh/DYo45eAslP2ZSl+tPswshv
HvECzJ2ZUGet13hFOMk8LvJSBZK/EJJsXPSRtZGjvyH7fa2e1sHXiNjzxfxbF0u/
RDAZAroBjTamAl2+2P5JIyU1N2xNZJ293/uvIStaniXMWNdvb1zI0og02Ko15jRl
AgHYgVqAj5JIHNeaytAN/j8ajELyPbWJaxSFDr9LyCWswTxqZzjgV0iszExpXicQ
9GbCfCBh9L3DxYofzme2harbd8uMF9m2EqHs937864VS+zU42vihu2kAOAOKPV4g
uJSMkqlqJux1+AzGzeOjtQhen/aYX6pXvidcE7P0oFlCJMqgrFc1dUPMuSz5IfTb
N8twGQgAhDBJpo1pChFfsD11+G3V0ntbpP0v/MRwLz1JS2edWzNOIwZcr8BF6zg/
vQriynxsT/rwviXxuOcDh/JOlktWPiMETJ0NRhV/V+xhupeVUgqm2+8O5rEk/6p3
voJvMTwJGt9t9zJd2+CtvBAKwLXdB5w7NemUDO860TFPe6atj0oJZ1cmynQwCYU6
cKbRb/AOCHwYxlJRMLntZqeZzRTpaJ0SxALnt+IaV6w+JvBVTJWsWC/PTGKlhjqM
p848fgsBGMwM7aZYVBW+GdzOzTn41ThQtdErWiA4Fyncs2FvxtMzJsYQxcwXEvPL
fvOQDiFS7gnA/AQVCzVs40DdRd2KPj1ju17AYXBY19TvxB6Ebl2XXR0aWQ+Xod/t
uFuI9zKOAcnymqJK0i0BpwZ4WCwv9h3QWIi+tsemSPkCb/7M65508WOyNgdRCRS2
AI/FOqf7eCoveqoDizR8mCaxDLUOU1Njh0Sp85JNux9uZuck8rTWJaJnnd2T/Fe3
Iu95CrHWXSB/Xjm0tTqZPVL+/Z3Rj+leLUWgEpyOlZ8HzaRRtfDM6S3MefmKjzAA
qtMaERYRD6pHdmkUkmbTeE0GPUxAIed0wfpqYqxkqI7a0e46AfaG6VlYVkeNrFXe
w8gdX/xkScrCFTyDYJg5/2t8GSxSBkpqdkX2mimeA4vcXnbqpFkPQ7sJS6JongEc
QY0Ynsa7wX9yVe8RxceqsaSDjbyPOkvb0Ui+2p98L8U781KXqnCQYKeRSeg4AeQZ
A/kaT8uHekh/PoXOo/aWL31iQ5OPdbGI6XaBHnZerEgOUHM9XDDk+y6uLvGDsp2v
xcNN3Rc3sb910uLVWy4kVnPZ8EEZo8Vv6u5VsBJllwDOV0Ti/X19Cg+r8/TFjU+o
a7e1hYqk4R0Etii+7PCKOQEM4GeD76GGP3ae03vMGHs7bqRCcxT2v3aD47Bjam5y
WDUfzlSPSgMneQZ74yOlo/iauSPMLjDo3PRJmYe4kTVvn+/KEBxFEnsbM/5bdqS0
IQqtX9KGXlXz7CpILAIXQMex67qstA4ac0PD66wWipan+d8+REFpVGLSVgSO5SYh
0kyyQko2nYGJmTCBpnkz4eBKS3bgkG64PeFpmjomGulo2kLXQrDuT1+c3snr0Go3
8HFed6UHJPlNfP/5nhx7Zau16ev/p1/oiYwsS2IONKvYrB7NsDDphbfQCvDMNmUH
8ZD7+w8gC3wUyoyIWbey4eeSWI584Mcq5vNaYZfSzcT6x28rJPZ3Mx5CjFP/vxJL
VSh87LTBm5/74lfvo+/N2fiwTDumlHZpBVf97DIzTJURUxtmsWTFDg18FEIdvvuv
RqEgUpImMUVTW7T3zcd7Nr6G/DXLfB7JXCC6bv2A6Rf2f6gTs+PcXoOJuh5fTdcX
aWCzGsDegsmnXucqKxwK3yMkznnhHUb+lN1qIo9nDYeTASC8Py2MhesGmRqBMElE
oJZnIXzCLPhqm07NJwDWTs2jk0xqcygDD38r3BcSL5e46pzPQ4hHI1Wgir0mFuK0
wH1QsH4EUIFY5AnKCgUEjFOdUhiJLjwG70qtogkPxPaO5McCJeZFMFVYOgLxsaBs
BGb+KSYDPaBUJl8ERAh4fUt+qh8tqcR6cdS0dgTvWnwN89jp5o+8Z0rOOskXpAQH
1dqnoOjm1A4mLCw+K+a0+MEMVmeSrL7DJw6yyAZxSe2HLk9rLKmRO+J3g66bsJ6c
H/UJszOYd1x/Nre6nnKWahlbR5H0FpaLkbjTMfJ6SE1EqFtO/FaXq81hkTTS+3t6
VeyaJAE5OQqpUDSqc2YEnXaJG9t7SQRP9QfzTE3MoPWIr3Wy/7TlktpB5ec+XuPE
g05RngXTSw3GV89jk2zVAXf0cZRFeGqlnhzkLoc5YDp97IeyWbRF1JvD126MtgE/
87qqB9YbVQr4wG6hN19OUX2rsekxNKhaNnmFnIap/iOEzbBgXCwASxtHEeGTyTed
pCxNP1tQKIeGeuu/Xpsh5w==
`pragma protect end_protected
