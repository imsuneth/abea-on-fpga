// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ec5Qj+I0m7T6b+WdYq8Lpr8xuUMIfkf4/9RTGouBSKDe0x0TovAtQg4LmTheHSIg
80zkSWoDFJ/Y/0DHM/ExHqVOirSYxeq4FWCNvCdIK98/ABF+hRld2PmWBY2L85ge
kjmZA06kBy+rncs+xUbRTqAoZXhwfAMYwKmUcRCcfF8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1456)
vns6Hq7I+4RqX2aSLpaa4ayu1NzeXAV6XSU6wLuMqu1rNNbVjvKfzMlZ/IgITcqj
gnj+ePSM348Wt14bO55Y7WvnvfQ+cYGBL37sbuEabtUYnLfwurd9u9fLcQSMiOy+
dHSyK+ba/twLkCozxG11EJ8I3ZmocGA4K7AE3PKsTgkGe1aPDVYcc47XL+roY/es
szI8gk75Kv3gP7IcNH5tXOY2tHZaBY+75Ex5Hcs4gMYisMgwzBn+l8aWbsVXtxg7
M2QcKLIkdrVAFCOYVbFbud1N+KEqwbqmYYSDn8r/kzSo3J095RFSaNHdkgsNSAyI
Ex9ZJFQgRGObShehRbxl8uzJ8PgieNvx8UT6PvtBnmeH2iF6lfXjzBFY1wDt30rN
GPpvJyXmA2q6RtKAkq8Agw1qmf294TYcQAeYco/g2XTQlESEuX4cFlJjTVWZ+Hwu
DMe1MY19U0MZ8MUprnY6X8THCKTe7HzNPYpEr8yqysqwnN60Ja0v39Dy283sgWTi
IRRBbNiSmH+bCOnYhqilRjJuiqKfwB1GkEACXAllI9I5fy/bw0/9tUNGtoDEDuB6
gJ9ueTBHTNJktlEoWHwI5i4x4Cow96lMn+imqzr39e6cu3p7Ib8H0mHlBkREhmj/
V/1IbW6IX3trWqbnMtcdXQmNva5wGKYDZp6GZUOdlnnQ2L0vRVzBuMEOFFLRseJI
Joys9kkuUqPcUoE4j32KXLl81A/ew6F4PQZVKGpQHuDLSvIepIsHQCPeETG+a9tF
vdnpNat/mj/lJ7VaMTvkwwKJ1rNd5l8p5Gsuqvsuwz1dcCfR1M3LvW7fFUJRXgn/
fOE6yKPl8ZuJRiA7Ox9G0ZVpLOliVPS+onxB4n3nHqAF2/2OEFt7/KjrmXluvDWZ
dA4uuW1N4Xncxo2pSZM9E7A0Cq1JE9zlqoMunKZopMoy0oc/prST12HKQCqb/Uz/
yK6Hyu7bNJh1p2ECpqp/XgqdLXIbyuX40Hse09lNViknecDsJtbp0HSOvZnDFVwh
FPve0y0JuVAFKyCCLZEAerhSwXH75JMjbhAiWIl0ieBLP9xYKSmwpZw9FOh15Bms
H+ab9dvTlCeAkt9Nu8h+4YaLbFRxFI+ZCNdaq1XlMd7I2mkOZSVnduk/cxRVblr/
LDmgKHzZULXOMslgASNq7//KMRzKQRVibaNQnjVZthKc0sPUbs576YgIzpiQEaXB
KM91cCepbxeKMREAHcPQvzDp76xleI2POJtvOcd1aqy4yeg3c8u4SguqUoPLPP5h
VI7VbioMM6ICPP+OY6GCrqeGMrVWyEGdBrKvDtF8JAMZT2AzGD/7tTesrnDCpTnt
Cbj8dUbL4yL01TFiHPdoK+BORbPHRuXmEw0GywG4WpPwKKo/x09QLO5RYshEZp1J
aNozp7ToBoWyXR0apdn0VEUiFviquuMnvoKb+M6zuXl3TU+CKO1U68v9HsK5I7EP
6OuSvMbZxbNMrERx2IIKq5dT0tSQo8UPWwKKMQa2YrLAu9fa4Sfrm6CGXe+2Jrxs
qnKkoZKqUricNcC8fr2We0I8WFCPVsgJDCeL2E8mWC3kkj7TjHIBdo1jEAq/ca/7
5IKbIdp6MurFMu2UQNmPd009O6SOfBNVQmzJCybza1HoIg+DXeq/kJpXP76ERS6t
4T0BoK+ebBk+7WN3Fbop9v1C6JKbqoErW2/q3g7V0LuTM8cHbrt+9OFw/H0yuwD6
zcPalvgszVfvq9BS7+IBdkYEoGKDJIe3wkABOopqv213QLCyRDhWTbgN2jTRzGWC
xJuKY21rA/CUS571T0OuBEYaqCykcryEcsRHK3qyh16KTlb/r4BT3Xz7y14QPZX5
Kx7t+BFLX1cn9rcoaa15sfn0YGw4RffCgTkaLWkwjFhJh8Nlv81kHqR9yzTU+J22
MdZXTjVtd6n2CWO0tCn4Wg==
`pragma protect end_protected
