// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:45 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E8FNHE3Ws4l+vlpgtyTmVG9DU6XfT1TJO8r0I+Q0SYCWs4HXhsl3uczlPGIaOEH4
FZ7OSP4UX8BzIilcNFJDdzVX+BdEL9pnolfs9AnDUamWGhBEci1D7lWi2aB3m2wh
aIOdPv9PavdSQCyG/NWpvyE9nKrWn/uVmzXdCHO5jkY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
4x7UJTKc5KYaTyJspbnehwnEHgvexfdJgUtexWgxEX/lagxkdEDxIxkVhE/04aDH
Auh4vG6eBLeQTmAABPFwRNGS1rBrIbC44bGzXmKWrwtuPu+AAqazdFaTOGIJzB2g
q0OkMxmkufIoOxHKWTeaqJb51u9ftaOgYNfYdDv4NkxjWkfXdkKxYZ9cHKOb8U8a
szyywU3kb+yU5pTb0LSO8QbWT5VdEAKhA9qajN2oersEQiqEt+lymv3fFFS2wLtZ
KnzzwKSGTppD+HyQbiG0+33zAG8DWXI0CMz7jEhbx4ruFyP5qZYgP5qJy3FnL81/
qCsqix+GnEdLUr0iiZX/Y+b7bzxtEWL2W3K5hJ2/pMhd3W6GHNqa3mJsNm1sUgeJ
zz9hKQ4hTVnN0icfrk6ZW3PczVm2UTG+4KLVQuIg91wiRx0snzwarNKp8QWByCBc
HtcDyZhfJMG91qqKAhu41xc5bKxjQ8+zOzEwB+9J81cRdK1TBGWmazfYfa9/6Tz9
Y6J+XO9DJ58TfNgkiSW/bT3f+mojAswYph1UrQPzpQVS/kYagX/UPPXF/zsF3Gof
QShnYJJp4vMURv6fJuEjnkMMrQKs0013Ccpb1Vck2QwBryOiz7UXmfQzZ7zoAsI7
7coYQXcI/yE4HiOtOlDXrljZ55yXhpKTTUZdrwoKuC2LLakbTWwUE9Vc7+o63M7h
+5WZPEpk09D0T9639dw6wHoI5v6fCSO0WduQys4qkUr40rd+8k613PiRzzjH2Rb9
nNal1hLQTGitja8z39fhBD4miUzC8NLIlSuGkcJ58XbHgkT28YYnmQWYajD7i2pk
U3DCZGYIwVZapQDmmYpjZNq2UoeB0j8APlaYTvP9vi7o/1lCFJZtX8fa4NsAa9CI
x5/2H4e+6AkUTMZXNaFt3UrkHnQyrSdpKGofG9JkfPmMkuYueklPFvCO6+/TSxiK
nzHtun17P+SJFuWWV5azxEmOluHMU6zIGc9iQCmzb/ZffJkdba+Tee/UB5wfKM1p
a81zhSB/aT0/c8ZTUv2X52fdOqUgdfRFO9HsCFawNLGsFQiBXKkW/+xSY35kElPM
mvr0NKfm//X6QMP9zVHW8R+NWdMx+nMYc6t+CI7fw2mmO7Mbn/zVwT4weFMJbSj+
C2Shex6ANyLNm0wR5hsgwR3rLlBme5B8sXbQVfBkZJQylq/wp5riRjc8mYhjVZtp
YQWU/Ywx3u1UGsMoco/L3j0eu89LbWOr/1Cmv/MTRQQ6tyM18Rzp7yelBSZX8I+C
jq/pII6j4pgq/si2TTv5cufuX1sfM3adYrWJco/uAbKSmKnn9vSTZn1xuygC7JeE
psAvirtvn+Lew4M2sMwJEoPJNMOM6w4UbGqjWmbX//kCP0gREUc6seY2/0GngE9r
ui69pkpMuVe1g2w0BnFWWFHLvj8FMMV6Q2wNDEnx/ubchLhXr3b+/phQD5hw0+I7
72giWE0UFjEfYhWmCsuUoBGYKoodAGplfaBzMA/Bl+J9hS1KlxktypvkOrwkSvl3
wjoMi7T4q5wNk9Q9lLJYdxO2utkuI4+WwfgcDEyKUsjnq0LBW9PTxwDlhYhLwLws
i1sVwKLNWYo/nACRUKlvBjusYHMjMduLHnbP7O4vwdU3cXMJZWqGm3G+iLlnYRdN
HQXcLEa9MUx2fCeD/innW4YeW3408ITLhHWeS4++8YiIavkGQkY7Mt5tngRfbJiY
S0K2GbmI2zvBBza8dRoTJYtbS6MlBVniFmJPbr6K4d+Bxemee5JqCjGjEH1MnuOu
AsTj2J7dS6dGfVbbZIs69H4md23GjRVmoB6tIkQN2yKHKsRsJ/s2HZWkNp3zYIbT
YsYJ4F1jz1md4sU7i/qKpRy3h1/rv0Qwco7vb54fGu6+BQSshS0LYN8pPwIwro9f
DkVrbUTdJwG0MyP4rx2p2JBVeScMFxrqNXnza23WbNosLZPBV23vVk28sWGRZvCb
xgK3U7qRWIV3LI2GoEOGFa9aYTGwIbARJs8iMsRDI6c3vPBkgTygM4ZQnu5xNTRa
Me0qo6ViieH9Ww7VYtArsstOEqnH2PrNA1lF1l3ipnCPKfsEdZlxwluxoB/nsFpS
MmZqZs9sZloCbq+JXWgTkFTDPQUfA9fsMVSD60jHrU9jbAevhQDzBHakKk/ZmqgP
MXCTRibLULPYL+HAku59ONSGO1ndyNTkzgTw9N90MgmBEuFKRG3jLRCRBejZts6m
3Ecmq0aJf/nZW5VfLAVpkNjeaFheyE8dQDTU9pjdtsh0yj1qN5cYCV7z9/R1egmB
tCvpsHeEZI8QZGLYBN+2b0PgMnm0N/+G8vqEJt/Dd6mDr02Qe3dhu4v3tEc+QIHw
KJmsZbX+McR+Uom0JBrx/oO9KTsWT3b/tVUCfwrypHHkWPchctiLniszUB5+OLMw
M4YRmQdFBLMWDIjm+VIwAnb2elJUwzaj+b6rCO++7LD7STPnejB2YDco+ih9sSEL
2VWCDQonUN3h/J80B01qAG29wCXH/s3TqDd+JFEYVuObZ78w9FD0loJuxhxJGfZY
JmtiWNGlf2EB2EedqlnzlsLbAdJVU/Fl29ENQ2leL0XH7/hxkLYDbqV0wpFqp4rj
6gmMOTS33QVxkYUDYsWY6QGCN+DqDS/WKgM+E5VB7hEK1Sphq0sm0lipKsxRn7Lk
YS5M8Bly5ccstC3hLvB9CYVAbTLzn68i7Sc7XVCKBDglgxEV8QnIz2VqYsGiuW5t
R3FcAWbmsVEzcaFaE1oBKcswKctSK0eFDgdFxr9y/CjzCNHbmkR3/DqKONIKkeYv
o7Cl1L9wuQgLxWKUBcrYu5btpg+wesyGSIC/QC4YXmCUso6zpapNhaIQpiu1Uc4n
q/IVXW4OFd3ga8I3uREnOaW+QsB372W2jFyLDRODyD0lL7xGqhZyy7yHXfweYiVg
D8uLDNCtrmtgClaffp0gSUB085kMyZJnP4zL/cV2RbkwBFKo4uJ6ZYQ8BP8l9tmx
QC6kPapoFa2XhMmgtWJRJPfefEo98oTxHPkeRBbsJgAM1mXeguzmN+CxSb+tXLaa
YrrBLa8bHOnjlEQiclIKC3nhLrTJ+zkfMOPLfVWcl22/6lHrvC+LaFmhciAQRJER
`pragma protect end_protected
