// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:35 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aL3yWROkj0S780N4riiheV0AMzoanEJ5ZZ7hWll4kUH1+XBhXGfBSbEIfGz30Pjz
ZnyALnqRK5Dx5ALPfe2X2+zBClGoU9xwP6XleVMzeeUJTuoxUcUktO3x1DpQA9u3
NyY5kSmh78hHIdUQecJH++jTwoU9sY+e5QkCPvF26nc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9024)
uU6+wGSKhidY+nZyS+1BE+2eoYG88UBHWHa9j5StZuKbUZNzy/PgZfoFrmjcle33
2R9mGAm1AfNybsYUD59VQcD6AuIL6/UjOUhLR6YUs9Pq5+Yihv6Y7OvISGxu5msz
XHdy7meqxNO9MG0XoRAh2SNNMiQWWeDOZ5X3k9DaKTRXPvia6ozaCXDUsgpVp1DP
wcV5w7pp/fRChn/HNo07wXbhAbBHq4sidAlZS/mK+7tq6vT1ZetThWz6jjXm40HG
OzBoDkOWenIMK70+YkqWey1XtFz53B6KuUkkqoSBn5jj9fm/zTIjfMEoNcSkXjeZ
Dm0QS/2R3814Q/kWhEp5G0YlU9T0X4aM6g48y5HCPRj3Gc9Mhu8qrm0dftKcZjqB
fsfthXcv1t8EHBs87z4kYwFzM6KkkyqKGdh5zBfXtvKUDHHqev93tktuoAyYPQQR
NRq+lCDxLCBBlIKg/sM2KTd+oB/fJwvGI+XrtbKDwAJ/VibueYur4ojBQEF9P6tf
hS5noXEdm0dAxZdy0b/yVkUrKMscODsal5+xhl2I2swCBHUV5aPYeBXLxszE5ZPt
7E3SNfboSVtbE2erPO5DYtedTU/msL+a4/2+T6RMT3xL2JrjvuN+ZNXl4GpjOxIK
NnMQYQ5H5fyQOGrWnvVVrOgclSyibQdjQMzcGHGE5REuLZv/oAH7p94fmvbY2qwP
MBb6DXohjyhcB1GGR/HWHkuyWEfKbV3p2QuWBMy4v6H3fve6n2hOaDr3/rUp6F/E
6pmmsmocWrWFuUOXUp99YtTvuHS7vsg5W/YBQ7zyfYKjxFuOGzUw4OKbKnp6lxCk
ZUh/0lYVuW2AlIj466978Rh1RgT/D6rfwxnsN1OeMdPyinbak1+4FVnF7l4r27q3
8rPVzV3ejQbYRFNXmUIybPKUo+XUvxHAfSwkSQofNJTUVg+V47T16PesZ6KWsjV+
EoW5lcIM0tl7TwTSR+KTtDb4aGw52Ulyuy1yejah50Tj/qytmPtOA4MOl8UCGtBh
dzTFstBGrno2olD0Pg+8LmQoWxUt+dcwK+Lpcy6YafRax6B2KyXV14em33T7UeDC
70ACAj7AlxMg2hhZLhsHrFd42YpyUY7+gTUml/AywiT3OeaHRyzsPRWVfUzwkwKW
QbVSLT+BV1sA+E+CDpES+ic0qgd189rk9Fb4IVe2zgqfZrflE13rUno9In4AFoSr
ULTKmMASTOIqRRggSmgPPNpNEwIJfKAUgb5THEVKsZZVs54fRbVdLDorZgZdhLYt
tVlxc3PXHe6BIvyl35W0R1E2s+mfCZNH+YuZK/lfiVZzr8rD6cji2tulYri80OFW
SRg6raKNJximmQ4s2MzEfY0OliGV3J2dylIRi46NJ00g7EY1SDJKmxrcRIUSilmP
U535wkWW/wCGEi2KBPedZVhHJm1glEoqf4R3E5vnUq12TnLmoKvV5mNCU9HvJnnU
tBkw3srKRWO7YDP7JlKxsBx0Yi5PN91ET7Fguigu5T4d4a5IH+WNV5+ZqgOU9Z3D
m+ypDSb/uAtxa3OcAckGtI7hXfJe2zbhcJ+exfx0Po75Ho0Sb6c99SYRg0NNcx+8
ws9qKfBV6AR+UCQKrJkT5HuAe1iA108REK+ycKH2nJ+Tu4wWVOb6t3k4vKtI8JaY
3eghTcejHcuWvKdlov6ydO17i58LCTjxYXxhdnfFSG9yzvXDZ+ljGtgxKbwHVHbG
kL60nTFVx8BERbA1QTWdN2Uf9e8nH+TdPGe0ni8o+y3apgrJqcTxKVZ7h9iGinX+
BsutDfvSXrQYgXPlV3TSC0fN1PzGZMOY/03FYmqCuwF/9IhM5C1KrxInt4+SwZHM
S9QDTKpVEIlE8KbwikAvFZWPbykIaW2zQb0aStJIQ78hAUE9B91+3rL+hZWiY+Qh
58ryOqrKXSFBmlUfLaiHKYjpPaKHOPr8vdF8Efbf69C0qouW6tt/dEPkFn27uUNH
OfJA95nVUlMLWRanYk5rBtKNt+q4CfLhaUwcAspdp9XtAW2CMsAXzkbGDAGLLZY0
77SK4MLnjfSy6zrCTy4IoEoVrjmbsqUiPafcPXZNsCnQQndMTszCYRDmAe8jgit1
GXDELQZdlZfHuJl2TYMkPFhFL7ctNZVO/wWNFpbvEocsxLOeiAcFIV+C1lzxW+iN
6zxvpMNrbpHxtQM9F8vdLFZbEONfFx9KLk4Ccqja12YR1Wrahk7muSwubEkfS709
3rHfWH+0YFLzxKIRyvGn+MDjJShQThHtmuHp9BonB3CijXJenZprwyvhZy/11O7A
Lk81C/BNK9XNUdO6M1mbDcWL9Qd/+uLILv8Ws91Gm9BGKcrp0dD03gvEUr5IK/TX
Zpvcp10L9V3pt5S8nVv30wQUhzn100gF+3c66pHGlWXqdA5HjTK1Qsdbl+jHylRj
/02WZJkwSM6GWcEoc3TKeG4De1LIw2+mMCKe8dpjQezhwod976mlawi0wN3WvZ7d
c1UZ/oKE6LVgtvpMzLeK3H1M5AZQ5aZI5UJoOw6T8Tkil0g4/ziV6Jw92M8xjnTI
i3qCAK+QrNkdYk7BcMjlETYPt/5NaSRHG60PJ0UJQOedeNcM7QxyYlx2sV3KGnA7
F6AdUgRleqlUui9/oG43FApBwyvB7FPXtx0GD2wxSXYwhUZlSOV5FNGw1FSKLimG
XXEjOtZWlWLMdKo59m4aJHLVe7tDvCrPD8LPDVwrIJfUQ5uCjIyGWcDqUth96wXV
yKMliPka/3DDzkCb8Fj0cVZuKMS80w4Pv+zX0T6XToZu9R+t2OUVCKR4ruVZ4FcB
tC2xGJMtw0bMJaaCu21O8vJ7jEhSuyPs5slJx9M4DLVfnHuXVrFPtATXb7dqzSfp
JDz8CD8KjEKV+eHMAPgSWJOb6Lxjs/VCjimden0KUweGPX8h6vvJWcHkxPCsXN5+
3j1xPEC+ZeaHVsMXQxEw+qtS1Yz5OakuSJw6VYy7tazTEP+loK7ik8wZGVF4bJeB
VAZi8g2n7dXEIbDNkvZ/+z7WBOHCXxSGOogYgM0Y90JgDB5y41aNQ28Wp+0FLn36
JlPhs+Wexd5SR8+73rf+HSVzngy9CFseyFtc7XYnVqvSUyE4vODqxN/X688sLlCJ
kONrIVZASOb+Oo4tLPCajS3gY9cDshARO0YTwYmi5jMrCLZBZhHUDBlVmrhQA4S4
WpU33AknVMuU+UVvq2bqhJgte8GEQ6VzzUKJW0U2df4PiDNt2XVFZLwtXgNRTCf+
Uxa1UiGGAlDXt4+96wTIHQJRFnz4EEWXH8KSVEhGCNrCeyXUvlG6f94cF+m2/jbM
kUT1pK78umMQW+V0YAJJaQbaDOyJS2aTJ3bTzY/T4kTChbKDoIB5LnVim6Gq9Qns
XBlwEi4kQbWyhX7Qtf31gVuLe3aHYzAoGtLg6T+kxQqeC8BXOfjw1Bw1Y51hrKJL
7xMcE9BD0MOoP/HsY3arznmYNq2uOkN2tX7HtcmNSajV8sImLzBdqWQh85JDgPdb
RJ/qbeEMB0ZK7yabr8HoOlQyT+0ajNNp/lZWnmmLpkqfluOS6CdqBsCiGmv2LAEc
xXe2vME8ab6OeRH1QbGDZOKbS8r0j9241++nm3tztkLvAO95fqMNhg/ibuOmKmqq
MOZs6AEK5bOSiRIGydffH5MspNY0sPqWaKK6m8jDTHK2BIktaKhGfUhNLX7n3EyF
eJQfKHL7e+ojkp0WwKN6Kpcjr4rb2OcZhdsF4blGbcIIksN3zdFuJjvTkULva38/
1Zipfj9kasi6ZrSSvqNwQUu0XgqpAERp3bEi111W/Fe8sqCu4qR6Dap0R9LLG4eU
kk4bpp3FEYUZh1MEX6mJmmNf3DqzXKPdvL7E96NGb7ozcfnFyrtFvGKRFivw/SuI
ONwISv0VCQ9CUOuNyeYf4Abl9Nr6ZSZNEWWk8jvwMSptXeatsdUWZF20k8ffdWYL
tAlPD7RO9/KaEsk+OAv2vLVH55vrGM7xVle1i7ccj0jFnvMVQnh2GNSm5p0TMI+0
Up9v7aAHE8OtRuRhOIKs4ex4CAQNBinXn7muDV8x+jcgzvQ37M0Ck6RfOOhHTaQR
SGvOJuyuMJNjBovL+SlCnXCITM4XOUYCrjZplFfeVg/P599YIrTGSkeHJiVurNFL
mvz6520QP/z+gGTThXJKuwcY9hO362TyhnMqBpwm5kw4h39pk3imgy9nzUsH8q43
VCq2gJ8MfaFc8sxPPp2ePHNsnXBYLSpyObkqaZDM/HqyYUStA98ZH4fazsFshRU2
th/s2Lrnil9V96nu9ZkAHWydE63fJgsHwW5OK64Ks8MBeWeLF0wi4fgK2lUTWjec
6ydwR4yHUb3uq+W8wOBdHpXJSfWuOY8ZJir+7hbZJkraXDd+BgAk4E/y7p5wJj/i
bUcANPxc9oMc5dUhmpfB6Fl2RI7eU9eCtkIwHennnL9tcJo/OyfB0kSIt2TJSAVI
rxTZ3M55+M457ESx32hq12tiTEAcsh57IIs+QFVralgUi8YC78d+TqGC/qHvBQ5t
M/E27a4XB0JuSy0C+GuwfOv6DXmHVRN1IsKYnGnLh6Oa/bEArPrKbeE2t/O+CwR+
5BIqPV8axPzZ3ABTna9CZuutejBZiw3dUw/V2ZkDb2Rh2R7VB7nEwGftXYSWlc5s
5AxxCQjSEZFwxz2kqQzSeK9EtEufWE5Cco1ez2qYuy9qjbQq1AV2NJie/e32JVOI
23eAEks9Q1UOyXjlYT+o464oOFioyiZuErlENnOHx3iPVOQoOoszi3zBCZKw2ARE
NuybEsjLmtHcflPseCmhEgD5jC1F4RDvHMPUeLZQlVWDz7CsQzMmpJYCRAQy4cHB
YkY504BppCHndBGBQwQtVxZ7hP+LmMJeOCyGlU0ED1MQLNylJ3jsC+bLjDYJRbRg
GZD0exC5BhQprM6in+z8dtixIF3+kk4B+GXNfgX2BeDYFEYCBtLxRr0U2uMvXecW
9UF3cls/xJ1EH1cZNbvxhb3yH0IOI3yinlqj92OxZ/PL9tlPxX+9FnIn3AhfxjEJ
XtgLH8EDref4kIQDMJy8OIpRFwIFxbKnaRIhEukh8XX+XYUyv9FW8jlMBaCJLgE0
VgqBkqXhMoNnA0R/+Qj1XJbkXhHsI0Ut242wljnFlEwK0CgbVIvHJNq14RQ/xKr3
OwkMX87NShL5VhTwkwO/KSQ99pZkwT99NWJl8b7UJEcfWB7yGVr5U3h6CeqyqZCz
Jeczi5Yr54pvCxlpZMFW3HnHZS2egY4PuX5YVYx28JISTHyZTVPsmqI6om+Y3nwm
U9/LSB6Xcf9FY374aC4lKvq5dZPBz0jiWNXxj3dLOOyzDtqDIjUQO/tYEeKtISMf
PBcrLzUjQ2zaTkhQgIJpm5qtQc8VX+EKXQ2HKu8E7QS7+opt4QDKHHYVyBRuAd5R
FJfeS8tkcjdhmWJXnXCXp4N/xRB015k0HsxA5X6ZO7+pNFZc45gXpo/7oJOilDyr
oSs6BtOWAW1Zn7Y3iIkVkeT4+m8PRSDDu1ZK8dtC+NMsV3xG6+h/0vQgqc1V923n
xjsQ2oe5m5yE9q/mey66NkUBV3UWorTErYeFt8wzW9zC2SOLst1Q1+51UQxWQFOe
Q7P7MMjXogGiZEsmoi+aiPG/vXHfeRgx8rdA3d5bPDosQqC9zcf7qc5ehc567EZC
GgE/spfHG/0wMQWL7MkzGsvrL2XhBkmjbtr86c5h4AODfJ8yNAW2apghc5trBkJb
l5xE5LLXD2L6C47xQgyJuJ1qMTMC9a+EnM8Uj7DZig7B1ZOJ/M9M6BOfeUB29X+I
W7/cA56mv1d1bE76x5XTHv/lejkEClTZ6R5Viz13KVhouu6IWQsrXjgz00rW3c7i
uvW3Y+g3Fmt3FRQDU2NJiuLcUJ5l6tpMYvQBRohzeg48Qtwa4zhevHyc1V/9/88L
nA70VZLS3v8k8pQxAdr5TgSHTy89vdqUQLlTnxAMf4r0L3UbzdK8k1zCwQ13oU37
bKEqvJyaDOBDnCKMrNcll67kMDdhstUsmEDpe0G9lkI9N6YcL6xu3A7t+dK8ElrR
iN/EFPDswzkoucEqNbhohAFgbHRXb37tntk9UrxSOYzQ+0bKkY5XuABx4ZqFSh/y
SsTImNWUjaZiahVx59EYqYSDClpU51dLswRNQY98Hxnp9jVO9gaVYdmBN0Yoxorx
tGMrDWu+pqb+BAaRvjmvYVQmyxkwzpUfjUBj1Mt7q1LyDcGxL8YaXEXik0ezOzpz
/uhCqo/l5oiG9aMH1+1yUAVFTpqU3+hKlfmpCryTNqByZ3qMtOM1IJ+PiitKDq2F
Uatz9J9Yh24loFubKEri0F08kZg4IPad71e2wqmSCfa8qTJVgS1XKbU/jFWlYpT5
ro7YolfJo+oIsv8KgOZyBEpTWH4Q8WrkpBTx+AMXMQGIAol2OG2D6pdNrIAzGu7q
8l39jceZqYAqkU/lSRpuguCA3mlyLRFbaeA8gfFhKrP7dRDtncLrBZAFZadSmKO0
OWgQmuL4ZW0XZYGnj+842RfmZ37eJae2T1BwMS7wnCXiw0bnuRgb7SNZYrzMNb6s
eSzw1JDKCS+e5Vp9Pm0EavyuZ4opV0xHfVKZhEpttT4oZPE6lme20R/lQ5wpo8+K
qg0MiPAXdW7uP6yFLeFr25DmSEKVCm+uHuM2WmhJ3QdY6AlyoTu/0W9MF1xPkzGy
FnrnI11MDb38fp0z/5y4BaecxSUauCI4LmPMox98GaIkLCaMGmiV95zXgulJqbyj
hIZunz0rWUVVqDwYenAwfUu42hmwi0q7vEk3GLVYQiWfc+5v22C9NWap/gbQKUTK
kwMhfaFpykIQTacdpNLVkd9ECANS/JtL83+VkLvo391pgtdjMPMafD57a2jIUDxW
1/R0IwKjvbZKxWXFRS15qK1AqzuWWOUFG1v1xynvIxjGeAHzDlOluHmmRbErgx1D
y6eQNjIjGcAgWgS9HLCS9WegXfbhZQmHHihkJcEeOADeGKq7ufmxUMiFPaYFB02/
BFRqKimKmxpqGonoJKnr4Sez7HesVM3bS+y+YU5C40gj/L9vZ5LeXV/AJfXBvlcA
Qzow0YiULkDmcAhgu330eF01PzEvyV3V9IoGjbvxeP2q0WL5y8zhBzAMjDUg27Fk
l0ZsRBm4ukDecm4QvIINxAx8zfoyaTrbPZDja9RRBkXdUfLY0y9us9zu+R/SJCr7
hy3ow5O26vip4M8L9wVZNcaTPZ6xBAboNhshOHjg9uBXhAbUSQqgf9mpUpiqhdmK
3dVTWzgOzFOxu53rhZO9uOm3CTVKrJRYlylqGhMY0TPqH+/euMPA82qfj1J6dEo5
aM4wrU7ZfI83b2Rx+hMUpsbKu3hWv6/wBDtxmN+5nYK0aBAiDUvgPrPcRNDLZv6j
FBxEpnru/uvKJ1GMXfVg0oQl3cLjF5B4dY/2VFdGAlagZVev0YVXsje79f7WfyiD
3esM4joju9DBC3BL8fQAdhds4J23py5CA/T+ajawhypdaXobAOu7s5bVBsKibwZ5
HMEf87iEcJ5rUCvd3TVNzifPLmGII0wPg/5UgpFIhXmGvKyStfgu5yMSQD5x3ZgX
PFbh3lrPeBxVcPLOXmSefB81Ts1tFtLSoZ+xuUBgYMB2qdJ2WR/UB6Zbt8MxWEL2
DhzDxTA2waT8syElQk6vS4bUris63q4JDnBiB+1P72A8cQhS8uM+8+q5Wp9bge5L
MXEz67oZZ8r7knlow1ymc3TrsBboPl//w6f2qiV6wPcYQOn/bUm6nPqJBnsyovl6
zjpRfyxV2Wog9rHLm/jbZc3O95OAZibbEYVOE2sMRr2w4QUu9wAF63KwbW5VUBzl
i8KsNyIMz8InzZni0swZax57zxZYNhS+n6/d0gCg3bkkpXwoAsiucPYhZ9Vf2ljs
u9b4S6Q9y1elJmD0zYtw1MLfZ1ANShUfzczrz96OGAk7ndkI1Az5KWULI9WL/Znp
KwKfTgfzHUX7AbZnyX5g5e+FxyX0T/XoC1MBPvtnA6GxkRKywEwOuCqndr/ZU1V4
DpgwqwymYd6XjkTeJ3UJGaV4o37BjvP2Zk11Zi2nhPLIxEhJvI68Qkdvt9RMeNvv
OpxC5w6Lrw+yHA9s+CHjIq1Mvi+OgOAO1mWGQ+38/WZ9IQSYX3P0B0otXBcO/BDY
8TOy82k0yPRWwKwToL6fgypUG16K8FUjaq3hmXRouVHJXzf70YOJY2NR0ePSp/hM
JsECnkRs0BItTkBkLNjgo6b3HvuL6uSMNlFM3PNbMaMZ4KDTLZb7N0CZM4Cp4wky
3TMlyyOMMCbDtUCl39XieCconWy7RiAcSl4f2kX9pPYZ6sB4vq4QaJWYjI6F0+Wv
LPLJDNgW8ejKvBiR49X715g8051TPuYYL/MBhUH3lrcolGidX87gbG7EoMOqd1oC
Q03wWLkJUJAmOGDZpDLMKfgXlo0zQBKviPCOumCszYsZKgRbtSs93S/qq/YmQasM
rkgzagqr+RbKWYAhi3DozWIQ1dJGeUFG0HEGk7i908XTnn1k79SLtlBWB6fRwdzv
A6AFLy0kch1cjk/yzdlXjTIMaiiFuq5M6HFVba7N7tPXvBPXI9ZH8UHPMLBIxmS0
/z3fuMoKBMn3PyqcVAniqfhu14xDuMkZzZ4rKAa4c7ADYVPV+sjWG4yj1IhFruMe
CbvPk51eH/P4lIIwNyuBzDM/wnVzrjcvg54tcDQDFJZOwrYP8W5EpMhhI+bO/aC4
UDY7FdTSjdxLMy5vs4orh7FSHHwD8nLR+ic8PFHbalopESap2Sq9S9PGneI1pw2f
mpeeuTZ0c3Dz0zu5XAMkgOEQT98cAPiuUq7pAmCqtkmfKXBFQ2XDE19flLTxk8Yq
DoCiEItLm4g/gemF6gZNOtAcSWalimbJgx+cOc/yholcm3jwX5a6QD78oB0zizuq
dkzw6VajLxc9OSOh7RNBkzGEStYb4cdYVkA4kNpYQiUdRAW5ZaHUm3aTWqLfDNiI
u+VfaEAOSL0OmIQ6RS30v3mM3EI/0IOGrPAlwhPX0opPn7CrNFdvCZ14jY9DOrTd
vLl5jDKYkoeWBB6dVrZPc5kosu4Rre6H4VPcP66q571DoywPZXGOZpK54rF58f+I
sEFlctedsV6D+BBQjlpIzBWR18jC7lBdBjzIDHzp2GvbnuLxxXZ70IwimUByMxHB
gDKGlnEZ+9AWLVnc2fwLw/eMGNwxyP2JjLeqEgTLEdYAp+1RKEAHg4oprY0Rb3WI
Q+qzoJMIMmk4pYVRTHPxgEfJxSc0i8hifDy3sPisKAH/TD6GROxEo6i7mvGSeEvF
N9KrNgy0R15zpXRu7L0hQapG3/9xiHxoQFOIrXhVUqOEf+bHMngMb9AtVnOCBZVD
hHECGNrewwRqI1vLjWIH8E3h1qWj6W8sZPe0f+M1sUKp8GZV7rFh4OykRgovOTcM
YfNbKYd3JYevuNnr9jngiDsVGDhuVZrLWLq5WMSjO4KynWDwlfpQM5QGXJ8YIrFM
45XAgO9lkt41T/qYnHYo4wcVXg0XvF8LmPBdVdaClXL+QWVTb6U4x+Qy0yooaGvx
rzbRK4xOVEWYm0FONVonCUW+lIwBQIP6hnuNId4jAB8UxDi2p1gjaa1c+X/H9uk3
SuO67CvBbEXO8zgJm+0C82cGrkinLXCQuz707/K4OwoiZejnq+p3p+U9Y17VDMQY
HMGKc4t+fg3lpzAJwzrHbpeZFqnDQxqYT7gd9Q1g68DrPIxPXxJ9R0KorLd0Mo1j
fkFGia4KAT/Dx8wsVXxKaUao1w9kWMPdU4a15IZFlDhuDfKSQzBBYKUnD1o3jiRK
8GQsnhjjD4pRGRHyOZM0Z44ACtpzNaZB+GgVv4cCx+srrk6s/XGLKcEuGG3xy7DV
Bp54bPJjgEyeRxcRQTm8BK3d0f6wNdJ19wBROg4kk/NJqffblYhJO7Pl81s1PzKA
7/oqEuaxXNXy2d645GSXiTvM20P5+EZeBjunPLrk8EIN7H8niaTYQri+JSmhFcaP
POAStLehWOXlC4564lOY5IDX6AZ8IfEKDhpkvfhwGI1hQkbpBiV1B89lE50u8cXo
EoSu1IRiEQM6zqteL52zrDOJ8RaKMAdeMSBAFr3fLLXZcIMeFdiRV3jznV7vglsZ
ThyucJs7oH9qN69wwnAVa81Di0VqShLF7Ay8eaWo+EtSp+RiuaT7MjWDekSbw83N
nLMwZ3n0n2jszUMIvAVG/fCmoWi0AUFjjzhp//scFjWG4UOhwxx94L3vOigt7Pie
S0BwXy8i0sGIH9szKgF6jDJJA0zOOd1Gpqei6tyFVCJWVxL+eM8IwA7xceVhff+P
m3lxreT8MFcH7II6caLUk2hTMT5cfDGAedf69XH6eW/Ej4mLjQ7TpkV8RqBzjHxf
SlndsGhZD8NNWoA41NKg10yrJfr65m070UxpiIzbWx3cXZZsV+aylPt8u/M8Izhb
muFhTOjOhYIFsV8MUZ9/5/mwzXzAfGQ1gLt2PaAVs+B7kcVHIZGSAafhwmdwd+Pd
PanCiFQsLB8GvCOU6A2xgvMx4J9gD1M27UPEG3C5SEpTqyPiYCdGNEczsgglDaLE
p2y8QFbeF+qb3H0CFYlE/+5f5PdtEU0o0DDSGoEHnmhMx7+iZwbjU5/h+VbsU+HN
aEYLX1TIix78aU0ZSvS56HUGTK1+Mx74TAqWZM5qiTqzAh3yr6KBQX1y727ml0l4
rS1BsLg7904n79PFmUIwrkMz6CHbHErSnR9C2BzYVf3RQ5JqbeHVgRo5ngqdnAj/
zS4I5CjnvY7+VseyLJDdSVlLc1KbIQofpT2lP9OntgSMTmSva7e85R/9nDaDbAQv
bYuYipHLobGxS59ftkwsJv3f1bBazbVqaV4FFGcBlB/nyy41n4jxqX3gxivU9SoF
jjp5Uk6LrTkVLa2iF6ATrVjQYO81AwXRoM5UjhJ7WM1WghZKobFXdmOYonkYl6HV
gaaz7+50uVmtZBHORfdKjK6GEZRiRLb06X91xsYi5ZKW9HvGcl2hZz4nhKRLgl+g
s25WsUpFkwPNMm9FQSUqDvyux5TpOA4YEm9uvTAr9G6Q6m6VlYrXs3QC99twIfqK
ZFWcaCtowqaf+c5b/ZuIOJcyIOcN3HJ6hAv6UWNZ6cEltpNRTWtJRqfEcwZYqYKV
hQtUuPuIYpIYPsL2ENz3mZvAWihos3uOxbInB9r3zsQmljX/95z11a6UG7D//sAU
VlfFWWVpOa7m9xdFrxUniy0QkunvN5ECn3AJvwpKCw6LGKkWtNFcgzbI/5UY0d6C
GrvCTct1xFlUS6L8z7dZSSv1IzOtjSDXiE6txWD2T22XduddSDKmtmZ7vAIBjVxc
l5MqE3boldAPdb7r+7Eg0+EPZKg6+tVHSRBaesr7RZ72BVP8JuIiqFC1n/Tlg8jJ
OH5/dOZmgX6oVG7eLRKw76NbvNCjC+iBwK5xVpEa7ldacjwiVi4LLe9ZaUGVcDt8
Q+k2FETtI7zLFwCe2v6q/zlXIvNXYJ1tIh7l465kvzXc7xfYau6Z6EHgo7H2SPDV
mgtg32lRy00hqzeRikoJYBVStElfc1KG+Ny4ZGxQ9GLKkNIabgtgOa6wWNA1biYM
S03uxE9XABqnZ0iHyc/ZpVGUH0vFiV2CQp304OVN81z9F08klFdEFQ4ugLko2wJL
38ntP/V1tmXwqenfKTaRJw+Xai7mvGlorfYqiJ0JjbL6Loe0q/TFETGg6emD4ZgC
YbmchYO9P2E1RR1aAgMtetIS2ko9BjSeOAIgNSVrPdMNqahls9OOTgW6CphC89y3
n5+WRZlrwbq4qtlHNPIIRZdBnqDtc8sRsqUIsm8APONJwjBiK8Bnr+bNSBlNzJll
Lr3rA6nZ7NyebJ6cc/0u6zzFKDW8MqzgZMTL/XKFo/BgDNAdzZplInXlGTarDdrm
bFMVsqwjYx4E/HB/pTQ1QsGQmU0wmit7De9ZH1Ui/toCk1MhQfjG152/x2lixsbo
`pragma protect end_protected
