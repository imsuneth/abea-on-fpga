// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:39 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EGn6OObO0p80eGbiGDHyC/ppZPbqmhW7POh93cfgEEQuco88mvkQ/DnT1/Xx8ktq
gwGZN3jjD795ggHpu2tNmG2k7xckFrp6RUg9Ty8EP+RSNa+nKqKA3TnFpAQO5k2I
0v2P3hTLSztcmJqLx5nXztQ/ji9ULZgB1DbmcB74FaA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5776)
e+dA2JAJHCOUmTjl2kfTFgScXFCoJhpQbx76BdrJqhIchz+TAsx1np/nlcCCT/m3
bHiQiDU0J8eNvps6f03ro97XZZxMuOTXv9qSQ3HY6gUwuNkLfDj858Mm9i+llK9q
xpVCoqfcFBnkvMyCdJDcwLCoAErbMoxa8k2BeyMN6HZ8BIpLCsclUs+Oxnzju0H0
NnPziUVMcu8dPunln9F3QiuU2fwDo2aPlYqYFDzItHU1DDTmAXD1uIiAqrHluy7S
YCtlDN8LHzkyJKvuipE9chVB+ZkwvUtITGNVSkZOLxT8h7xg2PVnV5MUPZ6zV45T
IPMgvFZLszzYffnbaz/dZZqYT+hIUPDALnBX3WjQmVbeu7rNzD2DYjaVUO2mv6ix
j+Rn6AAwa0tiMn78VnM+Z5sycwmKlmNw3XbppyQ8pY9jpprfM1vw/LnmfRYyKB2v
ocoCx/XAY7xIQofKnJqtpmigB9FLhX2ifRcd7Z41aKkAE3yzpG2R8Fc1e7LCcL3N
Pu0mX/NeZtWlIcTF2d6NNc8BBYeeahQwaibZVmK8hASQuonh0hSJhlpOMs4oCrBk
UhSMRDcJQD6/0xh1AaNxMwpWe0BpbsxMs+tq2gaxwyyJLtui8Olb8Dh1W98hj9Gi
cNgTvE6LeQw7HlEXH9+duzTXxKWsJXgoPCtOHbqq6cybBz9ICqw3IYpI6U8+FMAY
vHwcfeLF7QgM1ilmkbc3ytzlkHMrh1DAyuaAHQkI7D7A2UMaA0kVU+OG1EnSSBLb
DQS7wQyr+OtmbIg8rhXRuOjOHtv6mMJ5GGVGwuKbjZLsjUPgrTgSPNZySgr+T1i+
Q9oNNIxvRr9DPECg/XoOnbXlqiCXVDwQbEkjQo+HhH/WuFB3ewC0c/BLoZ3Fmv4J
AopbXjhoRKn18pPzjk4+2l/G4eF1OcKodvfkC1QATEOm5Ji/zJzH15ZJB4gNBdVi
ANN1eN4wqMQ7iiEYilW1zwSEr4ujpo0E1ZV5o18TzN8tY0lo51boehs6eVeCljeH
MUHCx99jK7RgxPNTudd0lhFqwggOcJ3DuIL/e/cIEyuah013OuaFUxA4FIyyD+nK
dYUpsV3QZBEbJmMRlrQOdu/IFjJpVlMwqiExUQFSg2fsQv6v8pOJH/vr4KmSsZZ/
1jjbTzrWpYOW2LvNb0ZdTgnPI6Jt03bQzNVeLGgUy9yzQFL6gf2DdBOg1u3QK1/m
1liUFkitSyF/e5wN9TjMjtsl0VCIiodQ9kPfEfRVKdGg6eIs500yCYnIF5STFN/e
Y5vjvToI9pKr1aN1JDfFWlGJj9WXED5cnllMo4KpDoIpET4no9T3AEfUWiJeLMbS
GPQPZ2kgiBtr2wzQyq0T7ZqCNtCcY01Mag79r4lYFzh+CKUVVBmZn+S5S8FeGeWy
mJ1n8HSZ5vPMU3tOLJwCKD58BdF8OQadtfFCfJN3vuzIPZOTmKfFhcDcPi+jT7kS
5Fh/S8NZuwtLM3zi5UXRGyur73mzbsomIdeNFZqC2R6/uUjea5dwwBUAzSvlP4N+
3zD/K9BImW08DJZAiMkLFIU/CLKZnteCZuxWsBJd36S7hG/7cLZbQdw+AQ4TS1u8
h1Cx4pwr2GhzhhBQqhhlgfuq2D5u3kptsapHuLFalvrXx1BGC69iNOoCJGRNUeLd
LKVJvlbBEYOsrYfeuQHoUeAH/kEeJURmQh64e4tG0kYbMuzT33n1zBORPaa/nVb5
FuY54eWKdKmk9iGhuv3clJz5NrDLg+CnZmWaRCOfp7lBiObUq3i62fk8eLuuhHw/
rHF1OhCCUR7HIXQQurQeUlU/DPMfEE5bGArE8gK8RzoukBOlFZ4tqKFham6jdbzM
fwJGGYhcm4wvEVDNA5cxiO31cQI+UuAonb3UbufpXs5iE/HyoPt8CYgZMR0c8rat
xVgA6YLoKagczSg/fibNDm89IImrA9Mlaz4HzGS8VsTlJLn6oT3vPc8AULif2bca
L/dBQbqsRmQgim/8ylImr66iotKoG39L7E2K3KAqlrSIHNxanxaOec1hFLENxjtu
/IwLq9QLlZ7osLem96QEcv9Wwjdi1uupZOR8k8MLZPsUVR/0d0eIRcCtFq67NLb3
CuXGd6D6A/HLd9GprVXOwxs2fHwNYu7qoELo+8tBZMGTojp3YZzPJS/paW9oEAS9
lDsr2db9BGuGQHlADIpU15XVaovRmmh9zhmoq5yGZmCPeHFWnPpBukQThbTiPnXm
shs5RxpXuLZ7hxdAC6MMWq61AXtlFsMybmRnpAZLeZW7hL+rDixh5Enj/7Fg6gMG
rRatuvHLjqRY93cuTSOr3tsjwCE3TfnazSbRdCqfyfjPtuCXpm1ZAVfn40XNkfYC
3Rssp72nw6rscH+LxASGUPLBrbO61DZZdP58NLABY+WEwZkXI3/+d9qxv5gCzYsA
ojGszfLjx8nu9CHPFyppX7rlbHhChvmBtLymKmv7jhDAbtSGu/rQXog5LJAa1OxB
ZMPZwGuq3QV87w8j492nNCNGwFSic214VkzZ04KdIVvC3HQnAl7Y/M7GElPraKqO
EOKk8uBRyj2Ha67DMKQO42LkpOVCP7iP8rHaT8UXC9FCxhHpowEsO7vlktb29XRO
eQeWIYfp8eVVRm/Ztl8fvfn9gFyL/Pq5N62doTtBGoRoBepelVbeYs15Hnm9OKDV
c4m/l9zG8FCtqg8y5zAWUQtOm+u2xrRBuwYd8r6jPY5rZIjy42pVi/7exmjafTwh
pWZTond9PHrf9fP+21XFnmSUz/7teyzrjOVQGX94FmA+i5/zDCoC5Lxgtb9hdVjC
ApQKKdSklO6eQIZZ2zWuJG7FVxRR8/Qmksz+v96IFve4BKkleUjzvyYFTizwC4c/
19uxYGdc1NHQIvRFvhsc7LIxmzOT9ZTP7710lUAhbZEyvRpkzs7n3MbXwFNCwpab
Tgy1pjuZQtaXIzGxl56tnRSSXFA81Y58Yii1T3EcplNBZg7jIZk2xSWspiKwpzE9
G67erhTxxvZDe1RqltVPDihA2l0glVaC2EaAI0YK0d3J2XuX6Lh/7qukYPN7IDVy
7+Z/O0XnC2rjM8mxeVxqTZ8F5mnoTXRwruPLFwCxlrJmTp9YSuf9bPp1MHtwUK4K
xJJPtT3StQ2LNY090fl13Cd4GRqYOX+24Y0jYLHQP96i8cGN25qfHsibHP2c9szS
M3AiFSS6Z+WGPKWOK/ZXqLUm011SSHqkJa408f6DgDEWQzKedwdUBHoaAbG8YUCD
0yEaYCibjWN8gUTdicc4h8UR8lGY4bjaj6St2m2pmn675QWptTOVbvAmLZvw2XXL
GprKJcLoXofiYp/5qdgUrphRq+auJB3T9EwyTy7ajqT24AuJuGWo0n7W/y2roUiP
RUsSmzdBOfgaUObY5fYfSkCPxh+DFav0FKN2reJtqRvinBR8F8nJRyUSsVptICae
F+YwGI/03Jnr6TdLEa5068refdg/HiWHjjGof5H++bZ6DpUOMrnyKz5fzDNsLcu5
fPE2vl0mTfuOLv2jItN+dy4jeSobz+c8hb6dWN9mdajieNRtJfxlb3YNydLnCLlR
7TrFSSIoTEs0HulcgG7WeqeFiLm2aYP6N8ROIFxDlKWT4PCmLCau/U+7nJg3JaRl
NUne+3LKQPY+JlfxEfEZD22+2J9S3T6+ujck+EM3rLsyFsR8BimKBvknLmeqnC24
BC/IY0eLHNc5h0AxLvkk26yAU3aA3TlDswBJ14gicNwN4e19djz5IxpPG6x036pr
TGhZd4/etc055W48OztBeg6Fp91W+HDZDnCGzZ/XJ+5EXyNU0WxO16FecKfV589o
VPYi5Bgk0OXL0Ydgeq2GeRX9UHjltHNdpSozGLH4usYZ3q33597+x4PJ55i5Jmi0
Ogzq0MhfCHzpuJa96MhJIjVqr/sUhkCK/Qc28KasZZ+mbLriN0JncSQL+UI3un1a
bR+bXpOFf6Iy6k4/D9BkLvJxac/c+g4L9768r7i+tkfij8kNH1ewlK2+Q9w11IUR
mtGHx021JepSo1brmi/KnExzYLk1xG43GyIl7i5QEJpLaWUGoAg9BJfduzgqeYNP
h7Sci+ydplnWFJch4p4iRaS2KI5Aki1Zhioo6gqC16zgYqSNrHWcOGh2tHNwMPgJ
UdWZsdhCJC5+trY9suEYl7xUFItiH3HdwWmktgRS+K1RhWFJT0abpfpPN1hLllEQ
cD98hPgxcAYglhu0adnxfTXna2yA1xQefWxiy7fzw0wIm4tLMH29dOoHqKcQkN3b
KjdasGybxtdn24E+CY33Zor5iv5dSlGwZmmgb2GVUBBaRfvan2aEdDOwbJAZ/9Yg
cp/+xKRsCtbLOmxNkOc7TR1x2hfTIAuqdeXqqs88/q/Wq+YMQRQnXN+HcFRUzRmD
dHpwZRcuLYmmV9YrztOYArheRR8HtRWweDZGsw4iHVR86+Yab1BVEhABtcTu3ZC/
NiviG7+wxDSIcRM4WfyM/3A/SAwkFT09IXNbND8HAZvs7SZL+nFmXgHVI6RlDqI8
MziUcxxvz7U0KBMdHvAzSfZ8chxqV15ywFtIWMlLttWwbNgBiSm3X0SVS2F0Ijkr
Ayyx7h0Eyjdf7WKKHRRE+9sJofJUy6MMBHuByxc05LsL2kcwv8cfV9G6AQ5fDUkm
gBMe+2iPrxEKsWBLQS2cLIBsf2CPYLvdkn94J0qgvTnds9rV40pgn4PxNXBbN3Bn
vP6O/aBOE915YpWWzOPx/UCs4nsXOLb87QyGi2cpdE8G+n/qcsCKwQrzxBYAqb51
+6XqM4qRbclUSVN+FoeoOtjJ9/FS9SeP8Njt3vosQkANVZRbJhnONE17UMWFMkOc
AjBRlTjixQMB7zreqjLPBDi893qla8JBjvungyb2tUXY/8sjQyFsD6vzXh9FOnB0
8aGEQecMY2q5c3/5gDzIT719ddPgIDBTDMttbQnAJO8J7uzA7ddvr9D6etqz31oR
yH3HW8nO1IOz+xpUtzuN9vRC1Tix4bQNimgJ9gyNbq+CMYfp+AXjOKonVh6cDAIm
Azb7uMCm62x4xfmfWE58ViGcZ50sHbsp3lhprMyQY6ghgvYWvIo7Ko+joasxzZRl
7ae7lrn0CbVGpLROojB7w7TbreujcXgkX7ipo6qcM4kyKw1A7eolQuKFJvmzBHXi
LQCA2FYyhbvBDAuJ0YoIUl0LDzSwt6U/sOjUKo72vPiL3R1Xp60jLAlWdql6AnKt
wXcSNDXcs2sK9RjHN1meSqO1vlw2kizURlIAJlB+RgB03a/Zvmp/VnSUC6JGztZY
2jzxk1TxDSnNAy4kgyC9RBb2Pro+Bf6AinW936U7GXWiLX1t0IjMifJDwlzyB45B
a9Fy+jFZPAwV3z1PIk4IlJuIQunSCxr31WxpUMgNfAL7r4YOl6dlhmxZQ3vK5/iZ
YTMCSwqKXSDc6ETnQ6ea6a93P7EASwV0Nfs5iZGCWE8Ax5UvaY8jDGVrEpMzRBLy
z7FVtiERi/p0AbrYZd58KQc2GTyGr0vBUvWLQdwvLEV7raAQIk/QZ1PRtSVbHfmL
T2IWQGeSFIOTQ+cvOYKQnGDYPuB9FI6b+oU323vF4I7RKQpPAK2L2mCx93Oxj+6Q
jkPcuQsiZ7OKodrmoTcnhCa15BsdhB0iEOZYd6dcd1hViqDFC9HYNCSIJ9CYJgIa
6aMEMh1bkV5pNh1TVuEX39Gwlv636cdxJB5y9fIXoq7GCyANa5v3JUyUBLWDVnUk
REKxcpWoO+eIkDvSR+rz12Gky5GjvFY/FKY3klrucVvIaRxnw3b1LqOEuPW2s6T1
HDY9qWR6tavikvUJjkWZKpeGRKr9AEvWKyJrcArJzT+F6bdiPPNCDcl5HSrrpq2s
7JOvP/akiTu/JmBW1zKmM9yy6rl7AiYYEeniO1AS6PxjZGF1RYeT9N7LE50NBNfR
sSijw8m1CUdGudfqDqtNdlXQUrndwEFzFh+HU0Jatyi/fHbDl80Xw3gNmQhTukOI
TDmKVjVpBry8ZGEfkSLfgTeb7Kh2RClyskg/nBIMYnGZqOA4snbTHNDcsdYtHthQ
r0JXmqe1UJEbTZiwGIvG0Cr0uylcVmMXN8pTdipHzPGUpt2Bklkt4VTpGVUpVJYX
CLSafNslazN1Z7SfL2qaXdb0x6dbJIEGdVEgoOCNYmg5NF9VVotVvSlF+gUs9UW6
nHZ8VMFqyZhZMEF/Cw2BRqkzifawA/j6sygMqRIXQjfzFkSryuM72879tfT31hpv
jAxy1M8h0vmxY0kOqxRLzQVngA2KMQSc9aHNgpTLICojWMdK1PeRIrapRlBIGlFX
gBa5L8IBsinoPmK1/mItescgFOoQheIAYolxQ2FilxYE/Ag72NEjxBByanjDLhXO
1kAsUaqgivN+ZjMO0AmTO2llUe7rEW3jT2614e0aVT2zcB8kdashNZaUbKebweD1
qtxEEnWZVQxZIdQNTs+wOOfRL+GJOsFcyu2BaMj6vhZeZTOM+xeGolzTTZw+IS/X
Y9hh6/SU0iSf8813bFMiVu3bs+kWe44BvdgZrZRZrNMrwccSo4SwJliwtifzG7yb
GrkQlVV0dDpwscgLgVOb/uxiBM3HU+DDyM5Pxxnlo4HJElKhSNWgHgBz/KsvwFq7
Bdenilhv/YZJaHwrU7tytq0vQR/e8AdieKyx91t8k7vEmA9iTjw25yUPFRLXQ4Lm
lD50NE3KWAwwn4+lRg2l72csUwDHoVCXA2SnVCB0NFhrDTIVrik5cFb/f/fh0aKn
kIEybR7FNsU3nRd/O1MWDbEF9q+6rozRYEk1t6xojVwasXE2XSHAHm2iK/9g5EVS
R9jLTBazmn1ElANAMEj36ZKUH7B0UiwQsumWQeKWhNt5lDbFRA9xUN+6Gqramwwk
uM7xqtzVUT+lpqh53dJreeOSgVv56mjm12FpdHgeILDh7rTUPieZwfnhY8qM+TyD
oY3TDEb2LThklBfrohI0RKjwATAwG2o7hGdD/TWV1pEJmnb0z7HpAjY+JE8295u6
tXfpDwEbdAvbWFOpDquixnjiX2f3JO56ktlQ/7pjkPqJzWgZ5i5AUGy4AzOVCbN8
bBh01ZtXQPeM1AKXgo8O1mR1P1zXeJuMSHSwT/JBPH8uMG1GAmNAq+dd6ErROR5i
KeZ2VUzvdCj1sLaKd/xcvgVInN9FfaUceFVUkPfWxSITEOxkZEWnvjg8cTM/272M
QzktsV9PwBlo5i7rTYFh6gu6u7SK9f1g16mgzVrpsGIghc9tKEYm41z/J1ha8mpE
GlAuyIfTmvKHj/5c/QBBFvjmO8gr8cTeqx8mmgghvdJzlCCPgCjgY/o0CB1Lwp5e
68nZ9SbFYiN0rG/3KoqOTEiiD9/R1Pgdwx6W4gzcarI+RTOpixfkpPWgi5hMGH+U
9RLxlOVb0IiQKne4W5B5bN4zz9Xg95rOuMkKLwSu0PJdlyUpVyQnalG2McoSu6Tb
b/CUkwNWWU3kr9ME5ZMu+OUtUuKD4q19efejwkBmzjBsyzHjtI4XZeUgI+3jWjMh
LO3igkOjlHjsKimkOEhD/XrrE8lZ6y3dElMOgXz6YZ5xsieRcNPRHsQ/kVbsXxcc
AK0TbPs4o9PD3hYxwIdKq379QIXMIe0wii2p3Ln7yyWrzDRf16wOggpWpnSL3Yi8
BlvYcNWKDtFntX6+VKtjpw==
`pragma protect end_protected
