// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:51 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CC2mAhBy6+wa9tErFftrov35h7ZqxH2A8tTT2jQyiS96b56UxX3vftfzsXcUbGfq
4Xsh44j7+Mu7kGqtnAFSeoKJ14Mxofx74BYqC3l8PFeF8kaWfdfl44pyegQEOHdt
UOPIGUe1m9eal0GKFLXLst0dtrM+Z9RIUiyqRkXEU90=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7072)
OOf/9IGP/C4tDyxLIyyAloBxd+NjDZI0oJH01iBpn9bVEjni4T8CghTOr8o9EWE0
TzYlKqugqCDcAM+dgr20vURzKMZIAM6cdUFvViBGmkovC1UlGwSEP4dzNOkgrUxi
gWOj/VlbANaOkMEyPAXnTaJepSFotyQUEovaZVbfVvCcGmYgxwHbBcdybq/ypeel
riynH1NA3l5d2sFV2jZIN/QlmOQqVrmBMDh/BzWBnM3/x0iee2YgL7QBAtVnwQRU
jqjHoTNyE9k5HP2wfWU8Eln0rx8P91ReWpwshNihhKSaPp7dmepbVbHhuk/1fkJP
Q6c3ZoY9fLyO2O7ioMhM015KZ12ClXCZsKDf1j6kszqEkTEF/N73AXC77epekNAH
ivPEqRxdpR0XJDtOkE4fJlKawX5PdM1pNWR8vTW3R1T8tUys4umcGgQp3RlcvhiJ
RtHO6RmY2339wgrI67PbGfNbW2gI+1xbNHz5I3tYsoIlaAgtOpHxHjTbOCyKbmEr
6lW6x99dFgO/2mFDoh+E2W9Q0Tb1zP+Ar58goj5/om4zWyQaYHR0DX0/AtCUK2Ep
yc90Z3eyDJeE+5z5deLyzZXXOTwNHChBENZnUo9V304TOIKfcafwa/H6H/33Cr9k
EClnckYC9bBLqHXrWqKDkby30pX3X8l8WwEJgqOkYJ5aE2AmRkbo7PTPfXTlhmGj
k3WPUP5y8JVeiKmLi8NWdfBN+sT2BZNOknPISWgivnFF6D0jMPSANvYe15V2ri6l
Q4vs3HnaIIUduwGl1VeK8oLTpmZW8gLImqBA2YZTMrHLJ45+lXoxed++1nW5SdkX
kme1Sxbz0xunZa33I6AKPrFD+l1scySwecVsTrXUH07grzeml7pO4GwNHyl9EErc
NMAC5x33+QZYIja/Bq52ibd9qOqqgDGZdYPXA1GiTLc9GROFU7BDf0/sw6GmKKwB
Bjzm8qFdWwHmRJkVehPGCQFcDQA4F1bU6Kvse8SBIWo8DKya61I05rOEnG4WaDZs
0M97tN5JHViXfG7ymgZ4pbViWLeRO/6L12yAVLwYO6G8Ij6nokwi8PCU7VKNN7Tf
IO9ZYCKo+BGFxmMJ2EoXCqZKXqhHx9aOLbIkoRSTbGQNm52KjhaHFdqLah3bm5q5
60nqZtvjyp3q69n9zSZ4bSkUqVKQwYHFlf7K9UpPSFohanG/8u2hHfRwpUmGklG1
pyuJEVDdZKcl4FBTLnTan86dT4r49RReV57uJTXQQn3CvVS+7cbUpik2bjV0dT8x
203A1AFXpsHhqjsHzg/qjHrb8kJKbzRz3d1JJmWl1Kklrc516w98Z/7N6DIacNOt
GFuavtcKMJaKP7FOupYXComIXObsMTwYvs5IVDvHPob2WIp88Wiz+QT1vkwgxb9Y
93wLuBc5q8QG2n+pMPyM45DSolInzc5ob5Awrh0qZcP2WocAJGQG9LR5HVSnhsTl
c2o09IOsjew6jGj5lkGDMxnKpFfm9zsEcWMK4HOVjhxc+fuZ878iipN7rEbzWhj1
3RFuTTgoUscSiJ8OtTLp7x1+zSDa3I2glj3tiz7zQ8uTILWpnPd78PDeNQLHfgMs
haMkekofRfAs+PV3ZO1xNRF5ThWnRod07+LdO3F4n1bQuReLuYZ3607OMNkEdDO9
yP5v+Q7qPpfEYWKVaEVs/460Kg7Q5Ak6OPbg5VcdJ2LXrmJoJx+UTSUgA/rYq02Z
X0h6GQ3pQVJEh2QVkr92Ezs5pLtMqe1HLpi5DIl1S7H6/fVDEbnOmHxoLdzaG4XW
Xjo4TVK7VwWvCD9dmpAJEIs7FqSm5xoYXXookLWAVZtoN3zksRgSU9yCiblAFhMt
DVbdsFwQ0Sy5BkvFtwX87H27KGlmlrlx3gSNCsaEejvhYqpC5UhGXOy7IOSniC+h
y3iwIRSYTyJejl/yaAwjAw95eKMHVe3kMDswb+dVYaB6wlPUgXBLv04HfqaxggZl
nmAWjC81V+TG1X3lsh4YPYK8sIJVVi1wrthjOUeB703+GBz1EYh1XKXSZ2kOrzzy
pP8rEW7leR+o0Xz3bII8xGwU9nVCE02b0myvy3ZenPCXRdChHmqy+7MZ48WTCv0a
BaCIi5tQ5PMN0P8v8AY0jMKp1/M6brR99Z/tHncFS+by/vLJ1VtdQQKVjjEzcv3n
6hKvBoHM+k8txGzQH56NTcUMiHCUDcmWaU8DZro5kmZSL9PXHqFVp8IHebFwl/aT
A78b2KLq3sU5JobJ0EOTyYlcAmAmPpZgdnit2lcqXf+rwI53NXOuL5DDlBp+ytY6
msz10hJ9vcJdRvC7Md/4m8Qy+x+IAWMpcoIav2QskGZq4IDgwJHO6M9qo3WYsMGE
7a/EBnLRZ6Gdb//RyPdTCEmRTEa6HJMZgWHfLdJvqFNL33gOdo7LCfayAzxD0aF2
WaGj81kuowCVP+81AYWLs9TFXJMobD52i7z/kdfoEaMHlo2LQ3rmx1RFhtssYrzT
8+Yc4XA2OzkWYymj/MmEw86fjD/DQUTLLXMTbFFLN2SLa+U1epQtwgumRL9cNk7G
7Pf2fKss+5f+VeT9RsPcqtWNp7VJurE/2oQav848Q4TuqbzI9u+dVpIZZ6BR30ck
dGVCYRBbHSPq9MWkwvu9nbcLwHYT6LcigVTCGLOB8R2MQZ8VYNzpL085UtU78EiW
O3etNfKPjv2NN4mAKZo5ND8FgZXnzxtmfu3VGe9X1FG3qzCw3LYmFxfkzlCgyBxd
5vDDKH0fU28MQkqJuHTfSE2uyRRHSPF7doBJ54wXN9ysxMyn39KVi7+wxpo/GBYi
EPgpVDknS1KByKJpJRIKnDAbdQFrnBOC7E3sl/+hUnbS999Wor8MoWAFPXchJXi1
6ivKcI4qP670RxMZkVRlmjOrAdzg6TN+u0+z6QSFXHfK4KjuS06b6rD2L8t9NPUj
mlO92hd1R0OdkHxzo7EgALg5HHEyn8jPQQnPm9NSMz8/kedr+XNUD4/jjYle3M2X
L0hpLQuB+s0qiWJjcw+3dwMyO3C3DtYnlvsv0oZlooGSQs8Of+PMaVMBOSc2T/3P
lC1Vjn0qLw0PGduVz6t/FW8av3iOqY38sx5rE1FxFMOkjvaAo0kvcgY3BHj15Vmn
75B1197c7xtMlWZtKhoCOjDvAhMd6P7Gq8Dyk0Ov3Q8KcQIxNovMAwsmxDWXEdX9
leZIkARSt3fetHwdDvlPFQYyg4sxgCMa52xUeTds+Q3Vpd2X/WvPzWCBJtHZJgKo
sOhz+pWSzEWVbyDjigdaPGQ8Ow/0mybh6v1g9cghjRK5ex7zQ1lgg8h2E1dEQ7P1
nWAfGrMJd4k4AKXmgSD/aCEhXM2X540z0M1p9J/M55YoNGlxy6+JkuF4YMWHIbIm
pFyYvLOgiD2fxIkmjhBi8jdeLyui4+8+KPqlvU+jewthPDE6zxmV+jRtnU5dU6Ci
GCfdpDysu4bEdX6lJ/elXM4lDwBCdb0KHDCyhyTWQYyVCxdi2Xqzmdi+kKz31IEf
0KwNWhpyHyw6X7b/3kMlW9zr53LZUrH/8eQFgYomNoFy0K/CdpKYrF8G65PeoNcR
4L9Fa4mRI1N5nIwxCfYmJl+VQOKtUs40FF2RPfn3uObyCbzR8DFxSJ6xFVpeTkh0
mntyXL3/6Q+DFuyvQ9cKzGe/IkAAonqV+1FUpdlXYh39Sh+sB82OGYz1rSHKNl5K
0xQnZ1GKMPFbZQ/rOrQLJXKdCf8ncJqyl9Bgy6X/fVbv6jo/UbHd0kVQugaeOy93
6rOd34GEMzt884S3HuGHkcnovkJMDWNo05DX+0cfUwhhiS3GmwNsOqEO9A2qwnLm
gj4UWAIEV9xj9awLdpALnVZFCS7fImSfRJQzj2SX1elSwLKBsR3AgKIgb+Y3GoI2
sFByDz9qVOLEMxhZ0LKtwrX6c1KWj+Ge0lJfIxRw24mAFh4jUnRyr6C2HTdfLcRr
TbdQKqDJQ/qHHILWwJcPxF8RI4le7U3xFhE6YBoaftKHJ9t49z0UFvpl8fch6TqU
c9JAPLPl4zEd25casZM/jI4esNM/tond1uN7Kqf2lV8TWZn+voIccxl79tgbxRv1
3XfUnQEd0isMIbvoOH0+TaXpe3TkoJjpDW4PvrEB+7Cf1MoSrJ+UhCnGGBjZxemv
uOUFQQTmFv2jHl9EazYjx79b9Gw+foKdpoUom8qSq5N3fGuXFkXPHFiyHPr4U4LR
ZQQ7Ykpr0Y1zJS3hYSWZGN5IHI87sBP9Q57iXAm0v515FPWjxm0lW03kCRO+b+rz
p8lQEdd+PJMH86J+6qm7nUTMz1GJp1rS6Z7O+J0kS23NLbssPZSMMEJWME8iM++K
fK3GdqQUeXzWe1ojAdXWJmUpDF7mdPgaS9rX8QdOzU8PZfa0On2TunK40NZihtkn
I22iDqhdkGCGV8/Hxza/chAMCaS7DRwZAk6+3zhAGkeu6TFLhJ+ncBYFbxWQK/UG
oGJ5VhQ3J1aTtLqZxSOrvRYl74/Ihe1e7SXsKHBcAv3CyQ7UejKADSueWk/RRzeM
jqvikIMTcofU6fiBaBYhnGMmLEOXFx4z3J6yhE1DMSpfmowGXYiDSX3I5ZDcJVDY
j0QuWvi2rXpiIc6v4o408frFzuj3t3gTA4hX5zhvtB5Vv3krl+r+8tmHK1LYgph9
6SCLJED1cxnUpIYOahRO7eGIcb9ga7gLJq2cf1+I7Aq8TCIv1hSp2UvuKl01GRNN
Eu0Os3fPaIwKjkmDOh1ddw2PnPdOdNAoNNBFyBS20xxc2pAsdcigzpT4ABqzR8gO
3RFvpsBkJP8x1GJ0Wg5iLMwFnttXWK+rPkDkqYHUDKnvHIbuEEv2vf+s7Ty/L2Z2
dRTjq+sY0e9gmcWV4eVYryY/QDPk3XJpDFgh5Mqqrm6SZ1URAyuzwmrHa691bHii
Y3z6sKtawDp0CbbIhusBoRr9QZ875XMyMVXx34RtflnjQANc/kSqfGIweyQg3le/
CFZrP7zWtKUjHHS9YcHIZUO7+foKl0hDxN7RRCDXxT39P0uyeFW/Yehg0HKHzC5U
3i5rABhku7r+iqQuUvazuO3hmgABXCbTkmDSK7ncQ1tIDZwnY5EIH6LViKLSvThY
Rd4qSLAUbFaA96pQQLgiu40WGqFF4gkD8uk+hBuM6wn01oMBlmcSqIPDynPhF+/y
R4s8dLQpaouayNat4G3O+gMmw4XF+xwKkKHvesoFy+0vNoT2NCtKylRm9C1rAJCB
Fw7niD/TFrdw6go+Vj5a0+A8nCMfMqgcHwlnVvoYMXRZdENx7z+0u0dI0jnoOAOj
V7+yamJPKPk8KUIazcU01uTTZyXRBjqtqqiQqfC1CW+woNp5q9beDbh7qNLMzqnd
renAKZSNRHcaQWB63pIl68vSRUuUKS3NoLaZeu7MtjUUR/yXVg4F1IGmmZ6d1dcx
oLm8M1RuQMFxNHZteH7ZsjgTEzOljP4Jqfz7LfpWm51kV3oeHSY6knqizlebRspQ
UnLlREqsncbXq3ia7k++OWtZ926r5wDky40QqjDQZW7RfNHa99wyj+SWHF3pzVyQ
iLQ5xHat5dBZsG/IWVYJNkjpHMTgypf1u8awuX7wHOokTAm1iStsiBhhpIOxJppu
PFTI2h2ikBXGICHraFxDtsWslRHl/4xNQ6lUGZ3zsG07qcx5LWCCMqzLDfSIwv9G
A1sg8T1Sj4AEYZwC7teljYxJpvWsCzDMFlW0MxbZnfu6oOsEJGdONFkZi8HYRNTX
PcT7k9LoeVHuTnupT4OLbdfkv8YWwfJTfPwztxJkBohjO+gHWdYnd9dy2jAD6TF9
Mv3blTbc7GLziupw4+U2L7uPBNdV61REsMQA3Ph/p3s4mu8XUZuw6PMmMNgaiOUi
vLIWNTKXw1PJgtu6w/6HVhXXctR4QY6sxfKMIMyfnwNd4gfpV4L/+/pDTBzueseM
6QWy3GNtV3SkeDvtiiq+Vpgg0/G1eBrlWoiWQ+Mg0+Xb/QKJb6VZfMeqqXhmUJWi
68GAl29JPgOhaJJTtVDzUM9MRsEkOCfkusUw+peurZL7r17A5RwJQA2uq6qcJzoa
PiqA7WInJQuaaE7Lt0ktjmvkqFCaSKmNovjU9yE5RwmNEqZQ6QVhnmFAh47RedSa
6pv1owKCv0LhJa1fRqCs+/8nH1VPA6Y2aPmpyWmBLqkhYQSyTxX/8AXMlocHuPLq
36NFKCND0JTpjha5sXqWurRT3OXv/MiDbfwWRN/inwURD+PzFUQcMMj/5Xpw73X9
BO4N3oJS74MUYCSwxXDk9XdvEmMDO95aXjRwMFMUJMRrFl27coj0GMXbmpJtnFLp
24M3o61F0RJMPDzcSiXImSSRy7APrF6IaUsGRKN63mW4efdsxTefWNPHK3uGv4Dk
h0snPo2pGOhBrmS44aKYybPmMKu5HEnuP2URPZ0MwXli9dN+/5xGCQaxvRbD+PZf
pLYuwRnNheQmNz6WNbKeyjvMgFkfoT+q/E0N302YNzWlz1N4Q+Ebl9JEJyVhsTlY
HfiS8aSCQ+6PBCfKA3NeGJIcH8qMqBxN8yj0buBk0OGQ61xGLDpNKrcHpL36MrZd
mYsBtjYHhDr9HkVVlp7QIcKykyuckTIrr78n/XPf/hGFhJkfQLgbmRFIaFKgScJE
Kh0k2ULIOEon0M8bIRcgV07NVzup3uimIGgQ43i8McD/Jy5gOOkINmCA5FyMXDE8
3LfbFz/42jgkijMqKStc1JGkJgiihpfOqnZqoCpKw6EwdTd67zLhBdYraNxEN2RE
pZfDN6HmH8bVpZFcbf1dgdEfghxryZVTzdVqVLamvh/pvfosSFvIQVXkKnZtABmQ
MlYcPRHptqg3U2fZjUCJokwR9G8c+HF3GiHPHmI0g/3v4bC34J9JsO/y3v0Dqkcd
Hn9hW4IuHgZViZzi57gfs7Dy1BJg0NeU8SLWXplwrdNTlHr6MBVByX36Pp3RI/Io
G2V3f63IBEPpDPtD8XrVyr8UypPM9qLnzc91MgeOYfl1u3GazT0OwSTpc+BDOHGc
63qBBQrSIUZk6k/Yjq+mQ2YGmgabTWggI1Ab9FcoBx0puEVP7t0+ITU3cdThMR/a
vMX7PqOBhIb/GcGfQwd0b6Wic7Wu0SPW78B9xpJQKm6VpG7UOhlnbWexwsWWQ1li
wPLNSKd2X3+i707YcDZIJyS6DLOSw09SpF8fxPeBXzxz2jz/YnGcWCHwFSV31VWJ
06onrJvjEIF1fpgzhwA6AjTWGKNi14tSdNgTajVUivSHPgmR4bGigNlGArZVELSd
iY8oo3rnIQ27jBCDI8QjJknVvU1LSWcuyvnF9LwRIV7YnbkFVHd5Emx48wc6qxkw
OrbQb8RF3JvVZqEHgmmhnh6O4Dzs3rGTQcKf9/QH22dBomEw/gQNx5V5guXqy1Kd
UdyCTF78vi8O4T40QrzbVMX5qUeRpvGJvYKdtUuYb+igAx5kpnlDS/IrN/543fte
0vEqdkLz4rZoiNx9792Fqz6L+884ODasKrExlBGqz8OyCSUobGMQLe+IV2X+rZpX
4bnXSoEFeSPWFCFgBBtEkAXiM/Vic7+xpTiZ29peRLBQ1KEtcveooZY1CjgC/BgR
iD0+8JcIfksCK310kVEKTuBCfa/7ismSoy/pOwHt48fKEuMKRznUc5wdPbME5Zds
kg81SqNYBTXX/Wcun4LkduWLelmtfasEe+TSUu6ahkJ6whWcd9eI3xH+qAz10ARl
ZHI3x+Ctb6el1uzKJ+ArSqlXEJ13GtniJZDeolJR+5TcA5AMEmTQ5+UgYSM0wLXO
AsR/z761NvqOndFBRJSF5OND4mJYBB/aDrz69MuzUuDQZ8/eB2METVrsIL2LFTbg
zx2zXFeSqk08JPCVSB+CW6MByTGZ+Fr7nAfPrLUuVypnPJU7f3vApCzCat1cohOB
b3kq7rDwKpWhjH8DQknn1DIsJBPZ3pzkMaL3pCBaOUi36osF1WcZCAXKzVbp/jl+
YdSPlRzxYY2+5zp4Jj++3/H954hsal6LeQVMTywq3eLT6C++EILhTt4GC5IcWkfs
yoAmj4bEkVB8pqQmDe/3BJfXfyqI427AnZJTOYn+tgDRpR+oq7zUFHnJh1SFtpUx
mgxfb1ZprP/xpougfBB+6EuECQPkJdjOAWGZoRF5e7u44oy0GSvDh02EoiwDGzSN
qaZ8o5k1WiOMrM29XosmVZWtgWLSsizAzW2CQETSTDxvxC9lXdaprAUs4eKmaAIT
1KvA99Rm26hRBUEVMxJwzsD6wxNwhkojmK6XaEMmJg7zbv4mMXuOT+jWQ/veTbr5
XH0ZQ7Gax9mE/9DgmuPd/9uNBSJAzMYZvabhuy0cbiIrca72i7dgOwzFzioaKRxt
nP0OzntrFBcyjqmtNfuoqLRoRwrwimgtIgA20vW+OqXtbLv+gMj+080zBE3ZsLqG
k+NHzdVBdN7xK71egfIY4024Ai6fy6RmDkk7ZINLmgQn9uZPOWv2fSI1VLI7B7gJ
SQh+oK6AHU7XCtE+fXCu+YkcpzCjALEJiAl+GRthNSHzbHbKDuEbSUqO/QwVRvWx
HOopNEBZDQqkjDSUPExHFXeV6qhXCPLLCHZN4Gn3pvUFSHVYenSdYDWkjDtZHjen
rK1xXNpEyQNvQ1aL7wCKTKVimyEAifep2uJgldFPvhLQLpHqYuCuHkcxlz8Q2Mck
GaODy6Ax9P1HRvr3zXpBHAXa+iOeG0zv0iELIiEbPhTWtOtQROFAITV4eyShrUu6
87+Ci3zImIsL8XgmfyQ9cna9wGixBLa2TP2b1KB3A2a4k7/TMbEiiJOaOiXs29KT
ahhmA51G6mH01dGN7RsvseRKEsHiex8vYsCeebHkJirh1rFtjUkvzCnroP7Ejp7S
2py/b4Oz9XYk4etxE85Nj3lPnEmXIc+kFyb6eGUQKabk8NEoP0ISV+g8c/L1dpi/
BR4I7Kx5Jb3EHyxoL5hCi6W7Mwj8+/lvZxsg0sZkkj5vLCZ50B0+YCUz5lyFMz5V
zAwyYJNT6mAtdZlE07AACgYPUEoByiGv20OsX5bQnmM/ASBe3nm52KqZ7eq+kXSg
GG1imXf2Hoa1FlkCaseQeMhp+yOon2cxB2v45AeWmPEdIJW6o4f5dcKcQvQXsO8w
/FuEkZbcr/riqdtWGw2dK6oj8RYKZhD2LtA4hn46dYDKGXJI/1rci5g0leF6vTIz
nTuipsnhf78iJWXOeGhoWX2//Wx95Rk7fJYuqsEXZiCqr6lpXeHwyam1OjrCE0ma
T+Z8ekYdrdwFHtOTuP6quQir+D3JFfqNMCmHqhaCyyZvezOsD/ozc8sUteTBaN05
GUzWO8YdzHH/LF221PL82RmdScCpbZo4rcOY60f2CVqfJzqVmarF7Nmt6HoX+w6z
xSGJ7XdrKyYKiyg2cqljEQ==
`pragma protect end_protected
