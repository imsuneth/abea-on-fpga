// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:42 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GDpT0ILFmW/TNKTfoac1vXdFnwjW+uekOGPKvAUrt/wwnAR9W6Kopq+QGtgOlnC9
CzwYtOcDxqAa1nQYYIh3wDh7W5quH47BpUknFrcNE7rS0vq5oOZGHzliS2tVRQLQ
hKPec0TwKxisFQ2SSGhpUhUygSQqVBYIG7UIbWMQhaE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5088)
IPWhVUqWIyPjrbFe7zA5XOkvXJYVOagkVStHgXB3gjPqbCQgQhKYFrA7wkwOd7B8
U9L22z29lQz7W1OHBhGceD6/zwIbE+/9PK7A5S1WHivOJyPXdXnDntK9zRIaFm37
BuSgtNzbCA/+BX5Xne+c/hm6zYCmo8m/AgFh4G5tZNdkaaq9tXfWyq3UK8pN6zGQ
7c5vUcb4/kCA3+ZkLJ4pBscSO+g2bi4wr6e/GlHmEUEQsQqTSPao5tdEJajCznNO
QdoK0FxQA2Ndz+W+TtCF1AJ97tojHvLTcEdv0AyKIgGDek8ii7u9CAEa/g1rbjcm
hZEpE64tF3DlGVtXGMz9Dr4sSa7TkdMq423aUjkPcDeG3s3mKIgIjmbFz6HLIt32
YDywQOFNNqC5p0kp74pX+IIwdgMB9IiVO1uU2R5QigL3eG16aZJtVpXyxzkU/0Mm
l5B5rpxynz4j6cGNCDz9RkDLM7WeSt+5cgscuY+IR738yg/BNbkH835xaEg4HusX
+y2LAFgLRk6jl9G7vloqT1dr4sHTbtXreSxpP7dY3sihSVNtX3fQE77Dih4pXF9/
22P7B7DtH+WrpSjTMMp9Oe/exIu9XMjzQJm8ZuBzzVQqEvMN/Sqft0viyepvJzkk
A4WMdZj+AFM2lCURt0t+2nc4XgcMSukkBREM1L+8Wfh3KNZUfI10HeK4i02OfV2B
i5wQ+0m+2MJdZGKzjelCGfHqOyLB5KDIMXd4gDviTLLSgFOl4UxP6cdQw4uNO7Pb
CB/qeCilyyLqQ0ryUa7XE7FJwGwAKhRjC3oHBdED2B3wVpgmJEMsdLyPLXpfSBaL
V4gY4h+VGRAhVaC6SP03Z/HRsRFOdWPWBN76JuHGDJ6OLU5FBaDgGGh+dVfJ7asL
/T8AdhRMkCrGtRz3RX5qdSDy44A19TVSQq20f7NAJP1NTNkgH3UhJgznes8tMZSi
WaXroztNAB45yrM0l6fmowP97o1lNMPd/tjsqEkv6NiBkHvAx2JauHf/b8VKiBpV
H3kSP3Uttf3y+691HsIdtdKrMfzEZpn+hu9bYfS99JmiJSsLsyx16rOX2evflPub
S1ndgU6Myv2fzRH7P05G/m6CxI4JMJN4Xl2Is6B6m6ot4jE2GaaHbozaHbsL8Bd+
Ga70HuP4QBTIfxMrcRE34G5RfR/r5opCQhgF2uwylwnt3kexUdTqQsNCe7TUg3kU
oi3HQdU2eZYY8hScvbyX2wZZaaSKNQW20STmLzFVQO+FSRRHexRFJcqhsaaEKwxr
qfyBEWEYsAmxrvbBZYT3SHmXqsH1Ch9ufcWzI7v6zEoP5ov3InTNZET/pBYNuuWm
54vCuy+f3fPXWxMMpESz+3h1Wo3pnnpFKxR5UfOjLLLaxgqjRgCTf96uzncFJ9aA
0zPaBR101CAMuepXtEY/oGNPixK0MfbtDLwBgx6AVGjMMw+/0OgAB7sI/xCm2uHD
MgdS4LCf50GPEDo9vGx0xKbDYcR/7+SMHuA1B4O8568RXsIEZ+LieL6xzleNgaVd
BZ9G3uOmqXxt/b5CfQqblqNVpDHQNWDb5ns1Wr+h3f/mQPAAlv2PwzxPmm2Cye4j
uRVEvTTCs9qOG8GHFk020lzB3bbXWFYtqHUTbsKq79ULC6D8YWxpYGTcX/77LAlX
pVCPrurvuD1pZ/DXdSjDlM7j9/XWcm2rUsILZy0p3H3+ZGPLl2KyoRTow4xcSL6J
IbmvvHUk3OOqeBG39Q1zx0mALxqIv0HjMgd3IEXx7uT9WaxtiD6xD40vtfLBTHag
+pdswXaKhslgAM9WZhcuTpYduv9u+YD1XqfX7gzTFJ23Tg5Cp1Z+w2iNK1jptufT
0mmujvkEhkcnkkblVRg3Ffl0iyeHXdfkx2Kl7DO5AvnMba0M1fSs3vuMWzGDcXz8
Yd/wlY8l+E4haQ8FE52R1aB20Wqgs3fylnVwSIXsVJtbow5VEXVd+B5SzAwvKDQy
QMlHCTfBLGFKNQGVV2hBvkR4qVaBPkZa+1wRZbiiC0kYXktLxAFtqz7mPPK0rfwi
8ZDUypIHnM2r1wLWUBUjLZeqWxD3TrrWqe/prib4BFJM6wj7l6fMG2e9/sVUxIXF
ulCSmzfHNBchXS1bJG0b/54T+tG3V4g5BqqdsKvcqODGZPfpMvflzFfKcqGrca+S
WieIRHmNo55HAOXIonrB0XlTPNg/Ojt9/YOoMqzuB9c8K8gDs8LwdOvs4s0bZpm2
DzuQssQ57UuqoqzE4+VHZgiOk3VCBbaJS1Kjk5j3F+u2sQEthdalNU811KY9txoy
PcYa3MSsjtBTebIbQyTwOCqSbo3o329brilzwbEjwR7kzSe7dlXqQ0oUkYzC5iLb
DIJkF0Tne1lF0GRAKKg/V1OGDWXgpje21s6gDLWNOb83qI7Dngm/AzXOLd6O7GKA
J+7XAnw2ZPw0RWZI872GXHRRfW4OG0vqPsvKS1fsyaNAhJ4d3zbReieklNfd8JXK
NyHIkQVwdeZQ2bEairJf3d8vVILv07V83X851W5UJ+e5BtOV6sYDp9o45JsEgAOY
RRcCSGCN8qggmlAlLEos0q1g7tobAf3XVTmw/fS8FImiHQTX8lP3Oo+l1rh0ZF2t
7OMAWOntkyV9uaJ+qHNmfiVxGOBMhnW4LkIojbr/NxY0g12rcxnJ1yuZRdasTCoi
jFUgTi0ud45wQOXCx2qRTUcdiahiRJ2VrV1vTlK0pUBgO9DEL2SL1mmWn4R79S/7
vL+aSvqahDZeDPSFJQM8X23BECrGSEznuo8ejsqEALqyaLDLpBevgvrIl3ufqHzj
xQk+XwwnEiBJlwNLdEFAboqBgjn0Ccv4Hr9DkQeFJDYlC5ruO+0v8zaCTPeHi5In
3QgDpS/jkR+jQMJK5V0viYhsw9dcK//rrdxZ6gBhH3AESYg2JB4ZzRydZ+uJHACG
IbWKw+mCP5SQgQ2oMx0BwZEAcnvY/8h8th4tlSVBixWiDOTKeUszTvQnOz6/OT8z
ijPodA3Abfe2M4umDkFZwDOR5Jt5ppDgmFWHv3bGwiw/24cT0KzqXD5uuuwCCiDD
cpNypBTDUzLtdYUnthZggAwXQegKK6YBftptPww80r5cLXrvuZ7operWlB8tk6bc
Bnk6Toda/JTGpw58ah2BNycQJcZDF869onajhUmjbgXQ8MHBGI5z41RLJYb9YDxY
Su/nzmnIRTgKnazCMBzpN4xd7sR4Z75C915DUTs14GrykCXDI/DVU/y6TBtNDJHM
ckLpyB9YTC2X71FgqCuwdtHwhup/Mhyl82PDm40N0XYzOygo+1xkpR3cOUP0vwdR
TBQ63UpYwu7XQl9UC1VNjj9TX1AYY00vXCQB8jKX3Pbxc7EbsN2KkKybZGEafMNm
Jy0rMJKlhxatM79nqbmlvpRjQtMg5rIKsjSdQ2CLby4i/5KkEM5gV7QynzwAVUsS
u3hNppb5v7/CGXj9TTie+6XlSGs5656D1nnIAjUtDWqOfPMg8WRM9q9zBf4FEE8E
xjC/7ZBes+Et1IC3ciIVMIlbiPfo6RV8Rn65eeycvjS897klzTSbewGgg7cink7D
QPgIuXcvBDd4d1OvV3qfQxxzBDxOKO14mxWid86WnkeLx2aylcDSDSVhA5qA+ab4
iNYLitl65B5W+rHCGUUpqrXFPTUIe/QlOhjB9KRyuVGcLN8EDnr/GzFdWDCY5WPa
abh/eGEQ5/v7KTXJ1L3jjqgulpP8h5Smaw/A3M/7hQn9FN+l8bgQDw2hievIj7fr
3vvX3Tupus2e+zEjX/iyi3u3DtE2D3Hbkkw66fhF8bEk8EVHSbtJaHKRwoVtleI7
6FTmO+q7iG9QKZiCdkOinPYrPZQEgwr4+wo2n1QIZ9EhC0cOAEGc4uUgfZEXj0j6
I6ng60pGy9XHjkR7jKZxKsH1l+T6vyTPSA6ipoYNxW1StmhEE9PfqqdpbehrctO3
g8D+zNaYWnax13qz1WPRWaujZQHY60G5t/ih/od+SVkUMCdMpde5YP16AOPvSAer
hKwUPQrMeFPdC20dQb+lQYhX/rm/j+vI8RFhdpBXnDinQWqrArz59F5NZeNwfjk4
QXnA4iOzqDZgI9FBvOnMyCfMTuvbMPPAFQZAL1GqpyzXI42ym/sgCLKwL1srM5u+
oxxjfhVK/V13N6DV+oKAJI89PDJnnzQZoXhYhpuONEUzWYRc2lvXsF5oBrk+t0Tw
L+QOqXghavBlkKyXt2VaaCx+f5Bv3ypX/9qnJBqCqnY9S21ctZDKO7R+4OqE+qKj
ac5pcwsSQzySZ2hQZo8bqvvj5wD6Hvw7kkOadXAw0ItWPBVDIm/S2bTZ8ig6sPad
bIFjfX3XdV1QXgDd0OKocsVM6W04w1wRutv9LzCJoa2QCg75wNZWIdFpL2s+Hemr
2Jx7DNtH5CAoJXtrJTPY4EZjc6hVuOhHUqYMBQMuTZsDyuk7owb6U8G7RMv4nVeo
6x2H9wrrAjaBsy5JuGC3SxbLUam+0IvcWJtaSIC+U/opZWldOmgLkr2oHRqaX2Rd
q+EpOOMJOmiq9SWweOer56iDPQLewnH7G7YE8XximBfQBoT/+mzVmZZXviIkwGH4
EUG1e29EtGTBE32yZw2Te2BRyIzZ4QjgueIgXwyNaMiEZoIzc2L8j52yf21jYyYF
7m3tQHo7UMaQemfddkRIcI2+jzalYZ9Xk8L+aQ6CUH9NHdtxvazICechK9XgMoYb
LkgXE1Qbnq0RHsaO6aPWhkkI05OQeKQ6kVAw7ql/B8QMIrDnIi5Z47fEGd4qufHa
SZbXHr/bopSoSpxp2/EsFtyCV1tlsRIazC7mgcf2L5VMnWmhwij4RNo1zdyGTxLE
JwAvovVdUEjJBThnPOXL1qU23u/Cidt4K4BsFi5n1D5W1Iti4l1kIFRvvu2nYFay
8EHWSMvPmLSznQW1aPvtpYaz/Fg6e0AsnsW4hq0d2VGfpmxklEQNHbo667F4w7bT
9cUoJ15asYJIacJQG30EdINXN9RL7sER9Gb41R19GssW6GTfVH1Dd/rLrLh0q1sk
7Sz/gEzjvcAEieCeya943hJ9ahpJ+NW0j7uCMiIblzI5tQKahtHOY4O0t2jO5znS
1BcsFN9+2Lb+WFD5yW90GPjDkOxkbDCJ+IiVF/2l5E0+M/V4DoG8JN4FcTqSqHAZ
qlrZTkuYJhZ1KjFhG7601Ju2TzLrTDscGubOwhC75Bt7H+mFJ+KW/GwuSNu8WnJU
yN2y7HqF4iGsW3L7oS2oVc4h0aPN/tFCGo5wpC43pFfy6ySchCD1j5XKUyMxD0sb
bMB4+CihIyMYb8rxTD9anzDDagn8u1hajZzXIV/WT8lMonMXFOaO0IxpqHuwLR44
KHGZzC2XmOa3+HwbaSVLmXBWWZZZA9gkD6zW6/+577lNQumoAx11MQiwfQw0QvyB
jIb3m22QIo7Fu+W2BK/VmzKbuLGW6K/GV3oNDREPwIhI+3hKufi+/LbKE+ELqGpQ
voeJ5quGGE9YY34v/2dAkhXcViRVuxZ2Mp4xFf75ORfo9UO5rJgvO3XdEOJC6Tx7
hRv/J4dkTKVbK4Kvh48y7zKfyaE55wgnhVaAzquPA37jGJ7PPwtDmVU0zAvsMtoF
nxH6weSO8WZuAOChIOu5FInjB6hJsED8uphMhie6GhjqDddVG+7u6iPNxtWZE3fb
o4VNJLVYu2mvyV0qr/nGtDPqFrPlBnCev42u8xNz4cUeKCLuGSywZN0oCpLzpWjL
rHjOAd86vNFzY3v8DF1Fm8dCKwrl6iXwi5vuoh8uTVn2gmPewpA67BOUOhYBk0kV
l5Db3gVMonk5cauhIm3Ho5+pkPe3wwm6uIb9ia7znO4W802YKe/F+CqbnUpj/jlZ
17Vc1LCHGjeBBCmIBNwheJxQVVcJV+8kLNNyMKXx5jCowg2iWbRBdfxs1PIqTkn5
RolEC22YFRwDiMxZhM5/nlz98/0F2/NBWwEucHZHO8Y726ZtE9ve0P3MTQTK3vQo
3lVvGuWIdAos1hlhl/gMugBVAplRZuTLdOpiYOCXCioC4JU4ORpmlKxd8EIuVnrm
0/QIaVlDjhki+tRpXG4UOygomKwE6IDnic30bKCFqge5rbTF5ULUGFFWG9keMo6R
pP26IiF8zHCs/hzycixdFvz2rZH94e7TMq16M5gT9BV4XTIAIv4rZ32HUop+DD0T
9TBi2dZXaEC3h6ukwbFB/ettaSsPka4LNkvLmK1ihXw0DTWgHRThbkjf9LXdVcMX
wF3o4/usBySYcMY1ctuTIVq2BX6nrEaxTWlByC1DbKpJTMz4nNhDqRgiNP25Clko
A7LJy4onozEO88ux+5VoXz1jWOhIHlaT/65jK/VerjYe8c9yAbZyxCdKV3EFsVDq
7rGMHscb2SzDcdbmCq+jz6Pz/5DlgAF0H5DzNex+C1WfeHAD937bqsEKf5f+bGSr
pR+JbyvsdVIGGpQaz3vtR5hhfhV/bIXPSQ/V10wU3L2fqsyX57r+uWvPD2GcYEv7
gbePdMb5xflYp5sMjYBT5kv/UACKRFM+SMCrca9IqCnHzPdDwaQtpRBjZPDP2Igy
dwI9POCM14AtiZ6vGYpNSAMNWNo8umhvEMfxXknsxKIyYszDgelDHRdPnAZndcTO
0/I3cgQeQQgegAJZVImiA3r4wjYlw59ou6PzK0GFzK/WRJ4lwAfUpNWpwxn7i0C2
qRlDkWa8/xA2E5vEzavfShfnzjPyNaIXsbV6+GNxlmFNkftLiWfp1aopQPeAszOs
`pragma protect end_protected
