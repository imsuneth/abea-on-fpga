// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:31 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eKGuk77PA7Phl3y6E0geVIeirxJPP2J+fsgQo5R6LbX4FLIw61d0E7RXxL6Ku9Yi
WcZZ4MMaeU2BSeGTueNvYM6s7aCm7jWCCWR+7vRv9eF6hkpYiM9wFKvD2bPtsCNq
rHuNhXlY/iVx8G+y7NCVkNG0j/8LvKlzWSa6136TWhk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
Gh82EOyQTOesFRB3NGv/dpQzIKqKNjmB1VXFUNeg6bitou/AVuZ5UJ6LHLnDM2yX
X+qU3IrWCqNL452plrG8+O+mItWdmbkR4HAcDEAVQBEk/k22hfArCkAZFqYP9oyl
QVgL/r57N4IHrpnjOu6KuX0UKOEzpKK357hviLy4g60CCwQ56N8LFZmaNXpzJUBL
XzNsgL0jN4GGBmzL1spzdF4b7KdS0jOsgpimDr+GLiLW43krIKxgQTWps+BSQMbQ
FTbzpD1wK6Fnihyd+joTyGiiiGM7y1LS+ucyLzoZmz1cEU5TWI2tqBt/bpop+pVI
oqk3xOf3G4UcBpWCJe5Q4v/4lCpal/Z05mPceNo3ifODdabaJmYjsi0Gc2icpnYY
TKmGOrDpRx8jIsajUvinYUnIqqhgo5L8a6rjgnTXEdGA8TaUTxmguzITuxcgUqaA
XdGNwjQqyJ7LOckoeNKKh/1DM1PthvRC8C3zAv+8TaOuNKB6P4iea5MUyCpvxPot
qx2F8xIMK0/ZE+dtnH4r5MUIWU6IBa38FJ8ln2y3kF2aadxfq3HIxPQpYXJkg4eY
utmk3P87soCSfWmfm+uHOCM1aOMwk6iaNfznzObjMXdipD7OoOGT4Y4mIdRxzHpx
oKBWSywH4E+ZONt15c6ANqb++kjIE3BcKtIPxBfPejLVXodUt2ZIHzzxLz/lxSpR
PJzEDMTO+mtT/9flW35LLA0j6scj9NqxH60I8efTRbBX8J4RBv1a3DUoxcIxOwy9
zupk1Z61BfkOQ433NtOPuoCNaimvCAH4ABlZhNs2AvbYRpOYn3VAQnx+V55TAJOi
S8j0Jlike3z7Htu+D3wjxgneo3kDZBxl94pZNwd34hnSH61imtzlVqV2nrk3zufX
VGSuX8Ni8mOl2ZKtI8xRPKEwi2HNkgrNn0/nWHRk9VhTT3NaLsKDXBPhfPJ0EkC+
WhKz0+k12LKPrfCgDM+cy/XeFJpcKuHvI36f5cywNyndKTvNRALiD5tWTiEoQryu
vcPnB+cTzXBkYemAz9IMWuohlLBMrVYB+5vV6ncMN+KT10BPbdIlnobSwjoocBQ+
vB60zxom2LRAOPQfkcPjJGypqaMrueWcK6eesaY0tNI4Z9JccuGQQqHFM75uXiNR
mK0+fMqkcbIRn5IHljzMbFGOYaQLK1phpTATiONICzLBSo6RWBBcBK/g+nQG9fnk
gtGnieEOU+JEY1C/k83iBmIy1lRxGSjOtk2a/pM3snsv6QJGN4PsLBdnFdXxjpdq
+4+W3fyOoFUx+Z6LGj9MVe00dHDcvQEo9fTVd02J+MUZY639EqxpuRhAin+hM5Tl
oQquNMaAF7z/H25JMCF/ySLVrGBQefQWxkT+XYOflQSeEFvdgGsqy3vm0pq1XdEQ
0BeMO8c2sjZA9YFYyeNOs9iKW8SUzwOYHiLEf50tXUNmlRDTu61qBijG6HN5a7GX
cemxsE/5fI/LpctAE/wa0778YzHGqYiQh3p+9KFW5wTpriDktIs3ur1q0onVVOF+
pnqatptW4oiYb2iswMuyISOnTVUCpgB95OZLmUzjqBzUbbhK5p5cNkxBL25GIkhV
qU8zBSfx/dQ8ZNtFNHOxgnNZ91YxHQ1L1udDAZgrxHreMNMa6E0a2N4KIeL/FZCu
W0EzSvFReNJRekIHa6us43F1lFVlnbLMOy37vJnOLczF1W2PUVJ70qoc4sugr7zs
NxYR/ZIuK+0mZ+6x0qzN91BKFUe/n39naD2XyoMQ/BOU2sEVwNSchhwGFTeMwd6a
vrH//1+c9vNXjNr0gcVYrwDbxkBUxb8KerQNXqesexyfv53Y7jq1VM7syZPK0oDH
o76cluZsBwkw/P+iXX2IuUcJTO4i9f1QdBbkdzwQdST1I5OmpKjGaJERF6KEDTQp
ZQeLOBup//DVHIkV5EKs1rvmnvlJqZfswbQlrhPeh8kbs/tP7r2npvgLj8pO3Yy+
TJx8m+HUW5jjEcwck284HWQrDH/LHROKBWB4yk+AsrIn8zrAoEM10jvqttPpekhT
jBuvCGKwRj5i/5UiuuwVsWEtsflerpNWqLtuhBDw8kHK6nrgOuuv+GyMRhtv/0r+
OvGYNjMPQQD6495Yqhl8Z2tIlz/tMjAj/nyomOygqfQvyxy3awj3W44/IcESFw4P
Csb7iX7oo6O2hJaX6OldNGXAlqJvnWClaro4Dc1Ag9PFNLf25VjayRrr/u+jyyoR
83GJ2kGzXpZNsBtanFgViptBKYEXLP7dPOM4rm0iDsq6uCmHFIJAhFG3HhEalLCO
+hatAqNkc2DXMSdBA4NQfau6PK9R2t4c0W8VmURaBfCavfdQcs0JKKXYmp1Cjn6b
+f+76QheSssMWgPaWdkDTlvUyf5hAbaXcZGf7WBVtEXVMakJRuuRyd98Av3ND7jG
C0uz7x/SO91NrWp3yWYs6v4cDCmCq1tABIqC1P1zVqr5X8QU4FBH6fcfCsBrT021
9rpsNu3c87PUIcl/0XlV0xGO2c8Q9y8CAJIK3A/zwVAZJdpmTWrWg/4Fto57/vb0
+RDzFPWwcXcOfZfVBSUCnHA5mncR+Xc+FatlqYYolUpTQkvWPKJfesyLD6KGDLgZ
V3jDun4F8GAwGFxqRvM+f5ypq4GvKG4YFAOYewvRzAV70oTYnxaOJlcwWzeqKDJH
2X4XPYwODkkkTUtY1WHQIFwsoWfHGEr99GE/TduNApzDSlZ4jLEy6Mzo8iU5aaBK
jXvzp/w9b0iXnDWRwvqKTF3vep4+uZ/CeZu+idpg7uAJXmOOHjTMO0YErC40yLV/
jjJ4Xl6P3BA9UhXoddBWFHo6gYAsBiyW78/KcaiTueEJ5BeA2MHSXi1rjAU4Au58
5QTIfuiw6gVnkA2PCgOvGIU925THVAfbfT402/IlMH2FI7EvMwT6nRRa9z54DGsY
ssv29Pdacu5rEsmKfQps+6vNDZTJIPpTcXrtC7Q2nGj7AVmxnEd5p87JmVIMbq2t
1TfbRmPoUKpMtSc1W20pXXeAhpXRrj2ZxWvFviJSuagwIADLP4zNBYLTXEq8K/4J
qwMre+p9dpazTHcA/Rp20IrhORLedaRFXoeUCXVwKoAaGB8Wx1vJbMCnhycNuAbD
EONXzyFUDYuDXh0uUv92a3jg/n4mHhlLPkrk/BXYeTY7ol9Bugduc3lVCzWg8i/N
CIm4KQ4NqfoK0JB4CCv+aY7GyFUfXFlv6pAoVPgb1y96FmPtSrT+bG1CPuxYxxwK
CIs65fYieTjFOTvjGlWPllth9AMDkpcZKAU3nBHHNckenCp+d7zQ2F0sdtaOZuaY
lFIe6hS5tO78bfsScHJft4yFbp7gsyVmwCYJWZvfBenSBX64ULVAkcQgpmX6hCXj
bkvlkvRWk3ByegUNmizclAip1M5sK4Ky+nwquB06Jjqay+i9eiv9Ok57AX1WUDm2
PFkdu3AaCeGmm1xvIlyhumRxNw8CqZt7UWiR/ELo9OwodOa+Ov/rYQodzygk8Vsf
v6nL7OgGS9EnVZBq3VIgyvhgnt0kHTz5ztLW7AXD5Q4kWmfYc1rei6mjsNwpcj6+
Jl06TmlgDcmdqtn+i2bMQXkGfnRTDgZOHoP3XlBrsy9UbWrRZeoM50eCasB62T4H
OTuTnSuFGhyRfI9Q7XO1DB6GvzeNutyAeiRH0FNeqwixNT7rwTuSv+pxvjYuykGq
JZ9pj4QI0Oc9zjhi15pnwZ+xUb7tbc+naXqL3BL/5mTvRl1UTdMzxKbFoJmARNf7
GeUi5ybvHZCO3xq8agLpRE0NH9Wniks0U9fUVgWDrB1b++P3/X4M0NP2VQn/+rqX
Xma2My2dfwqx6tLv0NBcD+yn9yhMtm64DDIld4WPluS82uANsdIFtSJxfRPwz/+1
hDu5VM2nZEJbBbjDl8v+qJeepXKY3xm2m+mcSCbmNuHnOP28jSITlrpn68qNIjrE
XUD2PTLdMLd1id+gEDt/OUKgkklHI2hyIg7ohBlDyEOoYXVmbIDUltH9X1QgvH6b
EorQFKxS8RA3GJNcxq6gn0VRTGwcLf7XtmuHpKX6AUc6tZohtlgsDGNglUChrDVp
xyrFSjPvBIZid15vpNEDYr3su1hkAmhAzOA+iCSNE5Zz+OVVr6PGFUs5zGro7eG/
UmcDEMFWg+O3V1sHMpjyg8jIiHxOMK5GO+FdL6jfeXE=
`pragma protect end_protected
