// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:46 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TysdcnAFPHvA0dqCnBaiCZKgNx0n/JVpNB1YoIods0mAGmHSEGo4X/xAyoG6nzHm
DFDt/RuWg9i2bPn0V9P8rDZitP7Ick/8PCGWUx3vQAXldOP/s7m0pQN9PZNCSrQ2
6UahzNwa0L8D05bZ0m7bcvjmyC4NftbQp2tWlQ4pvo0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43680)
1f/z2bkiPWKfFEKtaSootw/TmlT/jD6afMbCC1nrBAYRBzbcUa8q39dWZLUAOypd
kyLGUyYHch5W6eX2oJORspD9iA1ZBSQ1lhH1P8qB05IF1YZ5/0HE5YetOQxI6xpO
8YNkG8AYmlNMirpc1LtncEduAL/sczBS/5uKNN6tQuB8LfvyJJbffD1hm9Ap5x3X
o438JRSu0NBUrKdAX9OOd13SDSwzsN6exLjJ8sWItaEchj0MICoi8SU8VpQ99FSQ
wwSzI8hx4QDxcv4uuZ9VTvCsEsnohURlP9le6SBCSPQH43kHTKOOY+iNcDRwh6Gl
Ch/Noz4Xc4+6QlB7M2wA1BRHIfJKqVKeWCyzueuaB2+RPMBhWPfi5/qqFM8K0b1G
Q3V+8d2InSNniFV9vcldSUU1/YTFfwnUDYaGlg33zWso2fIqEA0qbrsSqCdC8Dhg
9QhGkga9LDHqQJ0Y3SuFRhCN+vpxOtmhknprl/TvLlM4J8kSbUKe7XpZDnH19ypi
9A6E/ozT2zf1l+2XcK7KPDIicb1rrSPV3jf/T8Moor8CsZamIlXctwsd00VLBpBP
xYAiv5b11zBn6RKkKf6u502Qmeg0KIF8T4ua6uK4+q83Rq41OyIh5heogyERS9oh
U9NsaMKwTxmCo0goFnuZcTMe1lzNSK2qQ+l+mJiku/dxV7kST/vZUNl+voTZET76
hLCStd4DEjoA/rC29fKOBmNKL20pADF0/aP0UFQbBs/4oZ9CA1231Ifid6+zMgJC
l6VrOxQlP1vQidSI2PoELIGZ+i0rOXTLUBKHIxhM4iAB5KAYS+io+IJ4eKXnl45d
BgOv1sEB2QhMLo8tYk031cnXsuEi45ekK5dsbzdsRLtPnruhSIStklWKBUpBp2QA
05Bq/rcPzZRgl+lvrJCt0c89Ziqt/QwfIlCrKlvCwwulaC/DYQsYbW+9dhSRYqsH
6zCcwwDg2AzwH8Vb88Gtq++XOoymcVeoWxW5YKzgykSRFdVMM6TcwcbvyLmsdcFq
HSA2JT+8lKau2Y+xLI9rLANBEw6I+4DrFz6YYKcuTZWMcWCPBToKyWoRQJU3QPCa
SbxKEwkertB8MCmFkBrisXEU4Iy2+OjG4QryHW0LyympBHk6MsGlxhiOpRl0kVLi
TVit8g59ax1IXAzE0UtqeUJ4WMdXy9KubeStb1STdr2hwZ+s3pDPSw9h4vMcP1dV
Whm2Y5GiBNRErPa7ukvOVswRd5aaeyidJk2yKMJhyrfyDaPek5Zm3yknxw/PwWjm
aAMuAIy9g8LeTqmQGuPqIf7GHBEofoYAcJU+4ISHN8lg5Uv9K29Rwh6mrobC0iKn
JbYUTUwBcQKlQa4QdfPjh/BShSZp18w3wpfxLUMmc8kcSOavJKD4Pubyyzxv8RHi
m6hWbdRSvpAVFMz8LeSeySGx+8Mutq/mRMmvPXm6wGTivwIN2Z7OKfcQ/s3C4pCa
UKeqTaR7yCWEH1FCKYIL3d3TqMgBXbGN9b36gAhL9QHSLIfUKKuUCAgxbp09dzlW
WEOwere0n/zZKZ88nhr6gzHd+6sjNNDB4Ujjq/loDbIwIWc6ZZ9en05b61AZqljB
RHzCYO4wCukFQbqxFiXAEPkeCEt0uPJzm5n0tRPnI7vdTVy4ftM6i5ajB0V5je+H
dOgtAfZaDbGaYW6pnw2k5JUyYaoCTF7p9Xc+0AwW7K6N9BaBOEZL4ICVkThK/9zc
8HRbPdg+nEfScYcQ5Z5N3MkqGPcUoM6sdKj0LH/iyaFQbyvSu7bhyHgfuf998UjZ
IKZNn4zU7E5YNKCeq6On3LIbIYrcbsOarQN4LAZt2oi+fgupCEZhTfTT/ULeJ38Z
rP6xo4PGUz7hXu27jUR7Cc/h6e7n3q+I1drdAEnyrEgrVlomk5GMbpkvRYyBc7Ps
QGpi55OlE4CifaMjz1+GtFrS1uckyASHQxFJnRJr9uVhNGiVeMDo4OZVtE/OMIUe
m1jOMko28fMXL0qyTYdzimxT5dGdQEJr1SHcsZYJKWpFOo/iUa3EQbcm7sl7pNLA
ct2l9hRuH8UMcQuOlRmgEeXmKH/ld1Ne5NT+QBKkXWw54hRKYwOZolV7doH04SPm
FSgsUcM7sOO20RFmZnXq6Cmf0d1NoWy8/C7ERXWmklvca2qs+xY7w2N16cbPehTP
7WMsIQtFIWY7SdNeO9JtqZvMymGBHaLuJVC5ls77BuoPDHzxTDT4HIQnn0+S8CTo
o+0ccz3Pw5z/HjkcIOSabsfpy5Z192sVdgG2e52+sZ13K0HpqK59qYHl9KsJCLjy
coDYmWxSUGf1oBxbONYdyYIJmB1cVLdG0JURahE/B6tPnyrep90KviEuAQb+x86e
cO4C4EeRfVnfanamb0geJ+1TG1xfs22qEkcm3mjzRZLdt5nyPwXUObXv09Z7YZYy
y9sCV7lyZgC3tlHR1ox57+EnSmVcXFYSqbcbNemjIoLErAArqeCy5dGJ8Odcz/EM
2c9P0MTNjsTz81WrdGSXmc4OzLNxuOHrndxjblqGrufamEtZD7X9dAuMH46mQwWF
ieV/pK3d6hGLJRAkwxnB0s+avEEqAOUAPsdMCnXEA/thL24p7UXrtDhEUF+XUXWd
KzUkOKMWUbIHHNSMqIwVWOpdkhG+vWJli0YipMEWbozKw/SZXT8B82/KH+QUzLce
4VkKSusI4VOGARJb2rSa3ha92r0a0D7OZMBI1TtrihCWWdd0ffQUZwOQfcHwR3Re
h8KzDTeog89iPxA2yVe4JUbFaiRYzvQuyL24UkUxGlHwQpw/Cqn038Wyc/QHQByR
7YU0KzX0eySIKFYqVam58QZ9D7qoPJmYjnoaiNiQnsAI05sZXcasi3DAdq/KT6Zn
2sleGjauHx49oInYu0z2nspxkFdtf5ocMCzkNW4PAJhPuCJJpjDCnDv13Tgy42ve
t8mLf82/Jtx+kjETm1ym9E0RwNVH6LQ/t4td+ZGNlibXXaP0xbjrxP8q6aqmkRuO
GelQRGCV0QR/fGXNt8OeiF3RZK1oP3lGkyLYF32Zya34qIYuoA/OGmfNFu8Ddp3h
fUchANVW5wcQXJQf7nLh1zIpUufocHxvvQ1lCuaBV/ejPOMcCrpA8EnNw8BvQNCO
+ZeC7yvKIwF7DiqGulVGI6wYfLAwYOxKwZ5n+914oPkBB6ogOs9sBFXXbHUZghiD
VoZI46tRGc76rrG5HEVNZsLSb1kZIqGaXy9T4/B+xI0BD5o1YX4vq0EvIYMP3SHE
qeGNNx3dfG+Y+b+aNsNLUogaE6TwlfPNH/ibVpLTQK5Di8Yh3VDw/cLCrpCrgQjE
J3zrZT5h21s8suAWQMfTAm0cenOm3FX+JyHw2xamdK0tlN1xdGxSpXq2Crsn8paM
I8bbp1zeI+BJdr2JVYAC9J2SxJQZhZiES4u1poNztTFxvcQPi8so8awWDUQvfBkj
/qurVDSCF8H4p0r7HzdJCkmenqH6jLzKQ5/082Xh5g3YqGfMYqjMS0emJ6cNpWrh
3snMgLq4mCdrT3S8MNWGoCnwQikM6UL1EpKZ0i7WlFMTWOTOSVt5Qniy6JsnhtWu
buPpsfewol4geV0S164B3yzizkDgUvEWt86+iUaBV4ibnD78SxIH1GG9M4QPjCpm
+pBnsNRs+RmLYgG8qI2hPFAapkw2S4iaIgOKh/7B7QpH3e55LozWxrCylGfLK7Kw
owzaooYBSZwkLXhPk38k4wZuXrd+3knzNt+5p7cYMeGCsTOPzXtH8ZD9HrtFmGFe
KXkimlavQEUyjdpY+I8Mm9Vdi0DBbsYAocCqI2AHpBq0ZfKcPqs/8KDnFNRE+DaW
M7Yl49t0gYjyd3kSgZuzjnD4wxdu99S2fWceE77adLwqJrVI49QmVttkW/L9FpZU
UoKvzbXU8nhYZuUCISaf6rWKjZ3YMfZIT7pZDrO+vtu//Jy/OrCZNwRXG2id17oE
rVovc+lSOkx5MnvGOevLDIvbnasquV8mdQvak95wJ6pSJyr0qha6+pR6lf2e7UEp
Ue/I9l0Rrwzrmm3C/AvIXfQstCS4lc67aPXG2v7k+1YCUdCLYBN125ixNQAfGo9h
3gvV2p/I/diZoGipNVrvPZ+GGkURbYscxUcJylzNDCk21Lp2wnEoUrcj/GpJ68Se
yDokkgyYtP/KbUwuypE0fRd2KQub60scwGb2IEGRUxfh9krjM39yya3xMpvdlDG+
n4DKi+OhHPAXt3ILSaTVUBTOiG1xCAwcRWG+G1iM1no5zvXY207OaZg3Zbt2iuUD
B+qna2Xq+4dUrYr1Mut7rN7pepeHHrc8WS/csptSftyURazhFUTBuT9Mg3aMlbiI
QGhX8Vk3GF0w+XoXAgy4YUOV7gApJm0Rr08V6lOcecY1rXuAo28IMhUDSXy6rzuJ
b1N/AEDgjd6LdTfJEkuQcJwrAfvC+Ozv35H89SVSdQB2eXI6H+FjDnojWjqXlZ2K
vuAeHhT0zS5g7jyElUoiUhqMcSUyRDc4QqukYXV/u2x+DfXw4ksBCIgXoUFt6IRd
OKaH3h21srQO9lfohQunp10vZSGtIJ7ysCxQ8jXb/U0QuJ9f8K7V3CqQOx3ZRBrj
GZphtyt5ASAMrFPGU4YZrY5cqy9P3Vv0Cad7NJkV6OQl+GAdGiSY6BRrXZ+41PmD
AjdMKhnX6McAuOsFevYvb/KX/wW3jFklaPTynpm8jdEbzqcSBm1YvU9FptKWhBn3
UfEtNDdTAik7+fFiTnvAWIoJkAdxvTb93OL2rZ/tn8UOTUtUIz+Vw0Nn/K1bdmAA
t711IBm2oZymlj+ATETzU403Ih8ZVABV7WDru2WLrzFSYtsURAU4RXo37PNFmzJ/
vxUcnbw6pjFF5UeXCRugXBGSkE/XSyuh2lzMtif+oZaQMebSc+o6HC4m2EzZxORt
EPsGeWDDp3giXZpVwMjS9qiprg258+F/LwqNNNSqgBCE2PTN1aEMXXsi34+Hw9EH
iP2r0BJT1JU7lAr6gcjml6QhikoDhjb9vCbJpuYvP7CylizAMNuvYSHZF6tNTDQQ
UAI82q2W8zo6LZ2O2ypHkoNzDytmiOS40yCuQOX8+5xQECjMbfdlAiQsNE9Q11xN
6UmLtVY5pAqf9zM6w5iAutOmloD7TRlbFQitLxvFwjVQ2hfDat8LlP/jGFgQG479
jhEhI+h+qmzCn4DIa4B3Y3eIrRe8sjEIY1j/iGCeIPhKOvrDoyxVWomq3JDT6zqQ
0KPJWHk/PV62vd6IuoLou0kcLBhKOKw2jmOXKSiFUD4SyZmQH98QrQ9yftil3arV
vs/rpSwOWcVnknKtmYKj25Hj9vI49/sK1kjWVlxlbpqkC991ueg4FbNAKRXi354x
Nx1QtxraEuUwI2G0EBQh+uDP31Paxts6Orq3pkOlG34EqJ42Ir7tJAl3GEtaUBiS
qsTi85kSQGyt4fqqj7FtjqMn0s4iSEqc4Bvuit6XIiu/fBQspEyOOgT52a4JpPE/
zmSkS8oO/EQ7p4/MxxLOWmbgn6fiYbAzhUhWDTlrlHUyjGXWfSjN3PBtBpkeSQRa
No7Il9oMcCyO47Qj4mv+V9g/3m0a65YzDOKWElUEWYRFefkBpgxDTOygfsZOcLwE
0Ns1sRb993LYZWhap3N5vE5hpFpCbPzcqkEPlu8L1LIYGhBFXl0rWgTkmnBt9ubQ
X4MtAhH6RGvM2p3ZlnS354Q33F1kYwjgCPs91MyJ+0iIFoJrEppZKIB8vXKtAph7
MwuLEG+ndGZ2mLA/1D5mRcivfA4OD3xdu2cWgVTHs4i00znthqYDLxvl65SrHzpW
JpZbsDYosr5H2nmQAzGDogYKC73OCkCXiyFtcseAmmi/XNV8b83vIm5qVxIOGJa5
EytZKDZWLBFboART/mijYejXEvAiUXVcMRE3kqfYbMJJ+Y1/5/BleWn2pAuQL/HL
yUqv4huQT+oUR86/j6ethmjkWmvRURCoh7xJ8KF+qEeX+yUq/gXpIO2nZi8pTai0
w1a8bk2y2pYN8kfqMg52zhxvyFbfjJswcKFtFH2hTm/FMDtJirm8jbIOolvZ9xy1
X5yH6usnAwcptyYKmGY+3/3RHdkJoj+XrWs/qWfL+F66ta7LxnarFiXI28sCZoXZ
E75bW+EGcE6mV0Mo8+B2FDmqQsrAuPIphYpCpS3KmMjyJbgK0YmSBqFt8Yq1n9sM
Koe2PDy6RZzpCbryGq4uv4yD+GFzkfmCLlAk6pC1IFXJLpINth1y6U8A1c7Cu4iX
dQZknNqv3kbiIepJg1SWTA/vP7htobC5RsZWcOTqRf1BD0HgI5LvXq5HF1EOxYW8
qiynp6mIef5ZYleiCanaUYUCzMHU9dZFPZD8PQYjilsFIGSR9IXDc93moAODXfSl
66Jg+eNnj5MO1cmDnaCe0sG0aP69+V8NmPcKbikhvoz8aJ4tjyg2mpEBL+9QYoXZ
7QLzm3J9R8QvRnz7nSfF8H5dJ0xqROF9D/15WKMP3KZin6ZTf3QzLdAKn4EwON0l
gVKeZg2kZ/+WiLdT3xn31gIMHVzt4x5A/37zz78C1DduTLT3lmM5Dj+MgGu/fZI6
CG1xyEdHX2p2kKDw6yT6sv+yqSzSRDOrQcHYGt6qTQND+c76umku+SBjv5rk2E5Z
94uT3PtRTF6Q97vBAjA2Q/h49oK/i2KpPLlTlgoyoCHOaVAAJJyZeScfKSpZHei3
jp8oPU58RjmfL7RLaZ7xbUfu2r+dxlYRuQqoBaGZmsPgXhbgLgdthX6jaMnH/eCA
EEbznPoKJtJXNMy2D9A1VKFXFXV3+dSDnL4Y2FUXtXtO1HtKK1DLUaPLGblfBfTd
11U04f6/nAQro4Oj2NDgvXliVXwws0A4Itj51g4Lsfekh+lOh4BPJb/5rds7YdJV
Z97vGM0UbyhHVprHdKXeIbUYaL4RlWqx08CJlWxmyyhotnKplOjdOXKGB94c4OCv
WaIl0xZxbcG08qSU8LnhCzCKCXWAZoFkUAwn8h7dYmrtm/pqUIGJcTJr1zy3q4vb
ntVYDSDWEiSN+FK3whnjeNn4r7CvmJBCN0wo4F4lt4aqJ4KjJbSz+DuqSG0FEP7l
sdy8eNMO93TIpxJfE/gArhwaCE7rrdB/F10nxZ30hoYCYJc5GT6j7blJNkIkKvgU
j/JJCDW/OE2kPoiFCQTS5QlYDt5VM38k0uNTlqJ5UBfCPT1jW2K1d5hVXCEfBdJo
gJPPcNYHV8kePXxDYeLvcz0nECqxTvfjf9zrkXSqetAumpzlCC0PNDRyZyvQaASk
eyMnVToHgG1CA61dUi07j3PdsOxei1XYq3UxSY5rMa5idEqR0Nm1V3GHWJFpbzHJ
e3bOut1CLEbIrfz5/48AHv83oius8r39koSuBCjk6AdQaexfJ73zwB/SUZRdr0SE
5AoCi0jLgMch88gPsJLVCQp0ggQMUcuLDlajkGqurOr0S6q5ay3ixpdMWveFQrEN
aD5KwehRIWY3BId5qds/hKm2g8dbzkF0NAUnt44XAGFBTSqV9EiRCZ3UcHaTadga
sSfnHSCeaNHh/3ggL4GT8I3B/Mcg4UEt3CZMQ2TdTVIPSkuQwhyxyo8kv1EF6odN
1mlI0Vb5GJOjCH3RIoFj+03jEqgY6OR4nbvYw1xLSx/uFIVOs0HpNzCvo61GFhZG
uslZhZbNwN1wt6HC5xqNYikydkTM5DDZwG2cWuY2XEppp57ROTiGFkyVIUQwOy0A
AUTPVDIr8lg95vfUoPetLJyQj+ADq3iU+0o7shi7jPEDTmhXzmQi/iz4lIT5elZb
IyAS0M/CJ31VO6KT7MtZjZgO0z2mzABItBGsOtlDpu/R1VySfVMF16+c7sH/Hcrn
gu0Ngc/xJufCi9E8rehRCjraTQRr1lSuii+hMmdXoaQz1pVl16Oe+YeQQ91sta3x
zAZZ0X9qzhTendygVmxlxe4EZ2bUwMO3ZwAuReiWLOJaRH/y5p9sDabTG+0SzYzS
8HXJt/BCR88fltY5hopWrnVgoG6AGAoTvms7pBUItwdPYZqOaQmUQAzJrx5AmrK+
Jgef40+dYGInZ89lCK5E/KIfxdxj5zCyLop01tRMp3AecbGuKVTHQOAOi9lmlROx
9V6SP79k7p0dWKKnPXTZMbOowUhV+sEH0ldkVpcRgQYB8cDF+WkCsqVIpxfnlE1H
4hRvEOhU9OjDGnIffZ6G1mNK+WToLWOubyzPJ/62d8cVnbc7QenYUMbVu0YBh/hX
ZtfohhX7XlWDLvZT3HjJpjVQsqOmFXsUtdsvxw1yzFFG+TD6Skht+Vp92G8xEio/
ZDtl9M6GUKWeQMCswZNG6+DnmSe03O7zWlEvbRMpR/luFg4MLQlZ3puGSvVh+Q5y
2pZUGMFygIHN9JPzB++s3/S7hDE/Rkcv7am1lPy7BMTXu6Yo6ZrLNmY9rEy4bge9
MpW70RWhehIUrFKdGM27DiisJcBWdwWv9fSfS51vZKCYCLQfFRdMYbOcLllfbycz
jqy7RF92HQ5gig7XAg6A3xoH3JtGLykbb7dYgrcoEv8p83BkSNFj4RD0pBMfg5Ct
IkaQ+SRn1lOxXrwpDCTZGpUG6q/dcb10Z8r6Gn4/7bCv96OBV+w46y5OKItyRMjE
oSh8njgFHMVTvhBsV4U/S43aIbH47b259gmKU529PEC2rgsDjbMgKUJ8RLWMb+Ro
pwk3FjzuYSc6DOCf+su8D7S6Qde0178B4ggl3KLCkx0bL8K/UX2uWGwMwuMgGpDD
vcQ/FVv8z3gVOYcxRQ0cE9c/Dqn1xhxdx4w3nBjqe05MiVzThYGllrW1ChfoZfTl
jlBJcL0P/2HCVFXi9gYKCP51gerk5/D4neCyQkWvA7wiA/VZSkRwOslFmxbhhAbJ
QIsvJdZvcU+Qd2FxXQs09g9xNEVafQ6vCunlRRlMF5lVhEjrxFBms6wDZGFTyWvc
W02sDcx+Qd8qsZ62x0G+ci3qH+OGO7czLNl/CovHTVutsJaOO7rfM6eEXK9asl0z
8+SXm1RaerDNUgr8Pc6pWDZrifX1uGKCl1byps8mp7VV5livJTLVGjxyVWRK0gbC
QaX83gm4EiiL7BQbHFZLcJS8Ofx+gXIDpzpaegbSxl8y/JX87srNIcPfB868WjWb
Ud9edecUG5ihCmlT8hj09lGtHm3ISNBeNT06EqsoKnOosCRkG0YC8NneOUsJBZqn
5FV9jx+3AaqO1R7S87+s/7oIcnBxPYCIFLAH2pYPpeURvD2CaB0XwfxqeOFSuZsD
1NjzhUmyoz0FJPh5vwgJBcuN3Mk7fDZSi25c44IdFA09MrItthGSTKk4wwhgJwwR
hMFMyoQG1Ix3VDPZ2/1glE1nAAoPN2WpaTAYTvYfv7ukr1hiUKz3EWUxg/dsvrGW
XPpmrSMVz/yH5vf10qcaM9RTmQjRTR22JaeTACg8rbIPJDPw8vsvb6w+iIeIM2Ti
OhLNR4v0FvMLpaA3Y7fwrQxH5vnu5txUXTuCfOkMk0tghhxR0AUo5BrA44pEPHoA
FJVc45ZfLUoCISolv361xroMO++S2O+eegyY9aIOUSXVCnnlbPdS1hEnFe/ujaJz
uui6QjaQ/wBTgGWlBI6oukQBFpo8rY9qw6OvBW/uk6lKk9YJXVNWkK765Yn1hiG0
3UA4YqeAYQpGWJH6SSqNkgJ99L/1h3HE8me7MUs2l2+fXpmhM6ixVMD1EzJIUtfB
SMfAPLx3ciAZ4gw+iM4vzHKDQxexsPs4V3Ep2qB28T5V4QfPBCpEuBXtyeBYq+9d
RiFUAh9Y4b6v1IkoUgV1NT5XxpPKV86IEBs8tH5t1nziWUvxqoNE4v+ON1BYnKz4
qNirXyb0PgdxVRB9RBoUmNki5esHBw76wFSU6fIdRuV4Neqf7fzKaHkeRkYEpgms
bzRIkHQ519LE5EpE30kCxIsoPhbw9q0KPzipfD//FrIIIkWoSZEWDiSeia4km+Iw
je4niryyf0AzST5QPMnDZClHb+VrNokYT3FteWSV2AhdgfA2+eiO2bJVppvieTVd
48ydg2CwMCDnD6CtSF8hsmfcPKw2kSBhfqR1sDLos96OnY/EBx7L+5kLZWam9SsS
Rrvo3qK2Cm/eoq+XCmuBGkhSbrbA/Lr47QTs0MYJpa7XVsn2X/Z5tMlWuf8Fkn6f
IvX6oCZD3x2kuJNa76gJhxsy8++RZNREpeUj8GFgZtcMwQVVtY7EkbqP91WYEfg5
T/+N4pDky8rUKyMa7wmILWNK7FELgr3mrmG9wfRlfteI6Eppb8oplmJI5a+u1qyW
DbzepkfkE4fEwZLyOiLoG9ZYB88i3jiXimhQaE370nbn2Rb8ckSlEmikgLP+EnDy
V4o35W+vOS54UAVCA9z5TPWEO1FCs44+Myswx8YkJVsNqqeunKcrDNAKbdaYOi6I
VRvjoMrIngk/A+AfUZadIMcBsuyh9gaBMb1Kg+HqwpnWEtAUDPgJysDJQhZZbsGG
jJm7XF7L9O8dYyz26qUgjdUomZIOYBJN1e72sbAHIN88GK8hcz/zMDydUwJTrwaW
UGuI13csSEr9sGTxNq22sXrm2Wqn2oU2vyFwK6amj3Ix//6NFId3/RtqQPEeqCT6
OTpMmXeWhRZFSlvHmrYqcQQQnGC3aD8IsQvqqltzpEijczACkhV16uCxIZAOR5i1
ToW0jcJdrxi655CmWPOdioF7HoEbO4mLsB7F/KK/FVCIPlDcjjqj04kPPLPwGPgz
drQvueWVDOLQEF7EdDkGqw1IesF+FFMV5J3OOv33xwAvzMHm/dx/2uSubH27yBk1
/DR13oNSNmk2sElpop1p5oMvj3YAatJTLSUN9t1H10Yjif+b+6MRznxYS2FCXqd0
ERmtHR0l8OHLNQsjx9hxf+GNO0VGpJGjS4Rpxrow1G9iQXEkFdnI+jmI5nZUcAIc
YZSs9Vyz5vlxyJCotzdM6v49+8+mEulu2ps68guRDE4a1VIWaKde23vZTJ4TCQz+
K1DyOBhsxot7k6HqNqUDKr3NuI1M4yzkKabiTY5pdOVegyPU+41WU3o9hv9LQI3y
Ijaa0PXPjjYgr3elaLyUlG/RDr+oO0jbgFBRnVK4VfQvH+tduID93zrLJuUIy7lV
D7vIFDotqIKBVdoTbv6w3np4YLBnZBwBH/YvAcgkQrHbTd/JwXHo1hmgjmWw/igA
NO4C9f29OUZmVtLearFoWxrB0D2OW22SRaA2CdGMH9vYMcV+aEBLaiFbyDKRaITR
VglXgrBQKR42LfmBPN6+Kxr0mSb1p7WH7HyHq7bLXyyOB7YrNgtYg6bvBPDcoQe+
1VkSJfc4W7Jbn/gvS9qMTtU4rq6mUgHLOfihOMmea7SUQs75Q7+/IGryDworYyxF
lIzVtkIvBJVt26BqyIy+rrO9uud81riyG3rBRWAVs2OFf9SIl6/i8LXts/r/zjbq
mtzNr7m29s/BFnyKwW6JSpdxBgNKAINlhBg77Q9YlHUIcZgVnUMpI04WPJjA5HiE
vO+K5Vm4Q/EIKJ+nS4dtAxVw/otXnnmAuoXqmmkkyq7bDfpoIdbBTELEfqOFKfoi
MAVzpSr9/S9ERLwDvFhpb4fHipFQ4ZVhFQ1IisWrotaTXkiB9In+CyHOAq2noFzB
isvkkSqUUHsUsodgm4MXgH7XjNdOwJFc7ttYRRspq/wzv4x70KWS8IM3ibBsQClR
wvMPmHrThHZcz3r/J+U/kKOMYNPMU29c4MinO6Gcow+IxAJWBgE/8mDnrh1mhNCk
8lpbYGzuhDgaKrWgeZRYRSIaAIAalGBs0Kfrn/K48j0z9hj7IxIVRd1JG0UqrLQh
kGQ4emRPUddftuBm6vXxgx3bNcQWbzkaLG++YvrjTpzlOmjOKUJBOLh8BoFyJ3n5
/3goXXS1bsaqAX0uBwiuP64o6M0UtVVa5MFg4sBmC2lBdbbZoF7/AMgkF0enxT/h
reip7pTJG2O5/uj1MQmCih+B8QEPYaPSHBJbxvjaOnL4DaKhXLcBAb34lvEsBYhx
IZd4+Ou+QOLioqm8dBVTA4dr8YvJqPwQUFgxcxCK0xLNxCECh4Od1JuNMmIViIS5
Q4AqiFi1Qi1NDuSUrebIGUj+EQIutNUigHRSGKnLfXuGYxrl1G5vmABUZg/qEQei
ftyS5RzBS1AAlVi1un9BD5Qf7xmDM92xXBYkVYC4T5F0/tlzkqI619V6usOP+grJ
gLtOGlFbKuuxBWO6FKTrAgM5ZmwQsd5w9zJ/6TUHu5wiSvVEEQ9NKG9lGB+CRrN2
kFzBcHqpYSEpIqhlWOyaymnul0Z32FeWelcV4Pe+a7VfW278P6BYXF8YlMmubgvn
MVK8PdgUXVXWRAA/p4MsQ5SXAKz0F1oIldJ0CIV+gkF5jl2B5QQL5FgVvN+3077Y
xGeDkKhAF1lC0Pe07sBMGK/evXM/OODi6yrT8ID2FDlddzdVHwk3y1rDV1myU9cU
P5b+oz2Z9sstG37kl2Rm4SczLYISFqbY0wPl0oAKbVXpfAnpSaue5IH05PjdhKJh
YmUzrlARDvLTdyUJFdT16kn5E4gNuVcxM4YAq513Q5Bb3ZPLcTzHSS6R1UK2XMDB
s3fQ5Ocx+37n50CdJ4x+yxjSA+sf/WVnP7pXxyP/KQ4wNmHXuB7GEXg3y4UOGDAA
OGSLdv3ncTUC0OAAnbUT/NiOt/zu6V0Mj79+OwmKbv+QIKppNK0WQtKZwwxolEqC
WlNdZFv7KEJ0y2j1RhxRJIgf/4tKMZVNKLWGPNY9ZPCHrOEvENGd1BkeX48ayq8S
MxcH4HLS9zGoG9eFvyQOf5PR3kivE1tUzxGqyaQDhLdJsuD+ds+lvJEVDt3cMkSu
umvAhPBIAj+Ts6NjBl+GvY83yD3ahr4sxEmwQIklsnWy72vjXENxYxiwGlFVCulz
oyoWC3beDfqabGepsZO6CFFb1WB/aNkq+opTupXu2POot7l/Q2vbZXaOb4P1KwNQ
otThlyqHLBUF5bV1lWQpNrm1PZrKDmFhD4UHyVEFs9fcGOM/ZqDHWYH1eq2lcpC8
/jDGCtMlKJ+m3jQxuui+Hi2QQdWQ8ojxPII/BceuF8snl7z5f96KaS6+dQs9lELX
P6TcLZJMZXzyJOMDgvJzlFrdHAXBvIxyOKEgfFiv2ZHPwYMMy5ch8SBi1NzmILE6
MNFxbTqm0cDmBNPkc6JLr9zQu9sBGT8USK+0Wp7XEgdu61yQxN/XVva2PhOyXLrm
vbWSQNUULHcgZFi8QTSeb5ph8YnWuOZXfD/n24M7qIfLt8qEhjWvSO1jxp4sbu/g
IwJG8GwyQb77Tz0ei5871vGkONBVTPkN+SIZ1cD5iDgYDXHojbykk+1AnNRfkxCq
dsYiRiOQLmAS5tiUIWm8WCRgPdzDZKmD8EIenLTtRo3RedOvsjY9rkaJ9rOszbmj
dSpUYM3uc+3euQeYBl2dUqYvfY1/g8tJVl3q/M/6apllyh2QgfhHpZLuQp1Ic6Ub
59U0BdoZUw1R0Ha2anQT96UqyGvspDdjpkCn/ObVdBAj+DXptpQWst89Bqk9inx3
v/GYrSBNsqHJoYM4PDz+ow6AK+fiW0izblj5itoJQ2IT9vi9+J0EbC2CTuL3bGr0
6oBqR8jVOBSRYVarqdTEm3zZ8ibNvZXIUpKlrEEzCXnAbdJjRc5Z5vPHIIzSMZYU
frtwmkm/6cQzjn+n2TXOD/0ethq3/fQkq07ryyTySxWLXkm09q8oo1OeDz/Gu4vn
rTyXKixzT7uEfai4kfEJpDd9q4BMgCIPJaAznTb+bTVv/CmLxLqJBYWcIxnJpHIO
6QDLmp5VVuggv8qg2zuOsEKPQ1nxfWpWhOoO4sD60/+NvvdZmB8hbCki7ap2RGHg
lT7QX4kqrP6noDK8+rXOhwKEmagC2IQVaf7Cg2d3UeeFeZll+ZXRUnL+3+tWlEDJ
OxIBy9np2euJJPXRAIEAwnahUSTxF6CzCV9kj9FAujLoKXoKdC7EjEXMn2LqSBAM
ah+eBTz8cNSVEIeG4CvqMK6q3YZWx4kmsO0xB9+foWA+ldMZfLb9UHFX5OzhTp0y
k4IB1ljAQPLzxtSTWF7maQI7xXg0gkQ86vKscLN6CC3ti6EwsXJ2UvRMsmXVuRru
CycCJDiHOMpFTrU0+DkjsnHt1wpd4kWGu5EKDpM8N1SSpKQ5Khw2V5w/lz19oOJQ
32u9rxWxKSesuRbJvUd5N3vH6tLRmNWVfB2MbnU7Oo7yJJ+yQdFT79s3KutwcuMm
GHAJRU2juyuD7gBRIviDu7JVV4qimtzy/2aqHOBVx6Dy1+mxYanW+QC64JE6MZJB
5/HDmLwpNqE8DsmdqmKqP/fQWN+eynho08uPV0a3ZGiCTSKAaqtlYy7Zt5wPo1N3
uyt+t8dlhzJRPJDVmxFN+YqOko9YtFLF73Yyu42O1qEILCHYxuPZ7KgNPSPhvXK1
bVYXhyYdjQJ7K4l3yNcm6OnIT+8TKpwbjl1Qy8tcCfGba2HNGijIjU087Kf82Sq2
93DLBge0dgQadO3caYbtVpGCQw103JccX3Khm+38AfeV9TTB3/vkcta1LHiyx721
YZpwQohpKQWHw5q+cnPfy4VszOwmiBw7V7Mb8tlzSGhYu+87F/LVPHrBFnpp46iO
PIJIVGJufHOkiT2+8i1fuaZYKhwvraN3JJ+3GGIjfZipzaSXek7znr8+Kh4G1XTU
HIh2LktDTsq8gM7TKovFwXAYy6+YdMLpWgRBBOiDLEYmoCbTSiv9URNNHtYgeL8h
vkwxVl3TLAqPK6V6z1tnyIOt+nDcUG1x5aAfgXfJJLumU4OfSXIkk1e2fBPYrQK4
vS279AUqrM4WLElBV9nEsNbDz1sAQzapQBtv6+p7/z/MmK5DdwZ1pwbT967lWmcc
aNlaFGgUnzkxVKwTmTdYbBoLun3xA3LrdOAC5e0JIkoyMoO9qWN2UdoI1yjUE3H2
KP5Qqf6Rhgnszu/pNkFc8gbt0UTOsVtVOtIR1Ju7Mi4IaPgTPVLdi+XP49RudoFe
XhkkRXwrZflWWpiy3bZQW/MjIiJ30C2HP/sXovyIUJMAmcECw3uL27H9APeuMgJu
Je9docQZCVxHUaJSzfH7WrYUiysMA51iE9zSmiaCsQS4O97UUA7oL/IS2OKmp/tJ
+1HddhKDBTFA+jej4uQKrBfFfJ5vkArGe18EG9Ukgwc845k5tIrSLRvuTdbVQxJL
kKpDYBvFbg+dQZ46D9aE0MbgVqUEEiZlKv1/9q4KSJvPPGxaRhcMkvDCscyAxGrd
hxLoY0LI//DaoIllSPXTxHqYdFFtWvEDQZL0u+JZAc13KLrtVaSXNCnS99K6XcfN
62EvaireceYXMl9G5ZxtFjryNfOXOowPcwoicesp/SUMO104BmBKa3AJz+3XyE/9
22OWMc+Mv74Laa0nas3yTzuVKVohbdFaEV+m0tRDKUd7U99YEzBnmmtr6WlE6wm1
xqbmr6f14Rc5qdV/GAOQg3KMrVRXQhTlu++Ob8iaCFonBS8KZCzunhfHga/fqiVa
4d0OHgy68sr9v0CCN6I1iMgoPnWfmg0mMoscskPf+TQ64u7FMVVEgA3xDMWF9UyQ
1s5dpVSR7f4FiqvvlS3EqYwKqw+4E3pxNLXlirpVmC9TAPCXvo9NJ2btOk95PSgk
0cs+7Qg6TnJzujP75mbOQ0ABeyKS6UmZ8Glyr0p/cM+sWtTdl4hVbt5WO9wk0FAK
aqn5aUJJq1wPsda3sZcpAodsGTIknMoPD0EDtnlsZZruBrAX1rl9buLgedu0pMtE
fcJ3S8yQAM3nCPerHQcCz4ky2OCAy1H59tyOixl+2aYoxDdID3UO2rn2+G0z2qY3
znk8pXRuFAe68Nt+HL+Va5ejfFqUTPGznFxkJ7ryiPUEamPjvJXyrV4iVaUtLL+9
GOohKr8BWN31cNx6n4WmEJ/uK3jZbTVJhBTH+dHyPSSHmBe0obUareiYzySxdrgt
e7d91sn7xhjDFKsbsVYBnTaglLWqRIyI1lX7ATbBwFbwhBPlhtkUCKCT9X6gc9M0
7bGHpP+UdmBJvoTZxM5NJeOFkVi/5ZK4uQRAVUP+jCcaNDzXPNBXZ7iuYXj1ByAg
nHXnk3ZJphSjSzm8vhOJ9idwz90ZeyO1ax1JI7qHfqgpYfwdqsyirRUeZIIzWcSu
KS0uV/HYZB9EUXxplL0xHymt9yUHg7lqRH/7tfBR8hFRAKk25I71UAJykn00Hd3Y
TTgEeZ7Q36x8HhFCmbvdomuNtSzpwY1DwIfR6uJFLako0AxAw0zuptUw6fZHUqZ/
Gzu8yIrHJdj+w9lZOOWJ/WOhkq1xe/RNb5ZNkQQy0vVUw9AsnYiCYWpWgLgodFVE
rz73YNajk8Fng0Zee6mtYnKWacgzlXluFheLGAIq2AAjMgJGYK3w6zG02xjPF790
j14VZ8ehvva2eVGweXQXsDsrrOWJpLMQnOq9MXDXPUi7Tx8rVeI0armTQey+Fhon
e8tq8UPf16NizX5iIqUc8K6TEoTQIui+gtmYNDu35+ewRFT5ti9VBv0q0tlBZEsL
TXk+HKh13cfAjQXebjUu7JZ7ysHhcaVLMotCM8JXlHEytRKfATPgqDLASbYADKyR
MuwTgzoypghXENEGp4O2axYucQmciN4rlppcagUsL7rsdjha5IO/iMsrsTUUEzll
uO0O2YkKfNJVEfAazk80ApBF3/DD5m4iZdmuJfDWlE0mG7sV7v2k3uLeUxpuM8Fz
8aGSqSGxt+Ol+duMs3R/0hkW8wD8hAeFfqThk+0hbCRfxfMNN9rg8kwbpDR6tYYB
uyt9nEeGqpxGA8ELqikjCSGfOdRMyAweSxYPZObYv38jDvWLop70JAnbbLqz7ssz
wh+IgPTBY5+YzDyZhmyIDUISwC09+Pf3sIpEweoMPssKDqr+q4EoRAMjlNAh+ABP
TFOQUGoWaHI+gxZns5IZ7XCDcfNrIgKEZJ30XofusFZLgiJabY5Mu26AXSrPBif3
jMSnsQfT/b1SAcL2Pqf4CBTnyhWOOsMOtcW4opSQKf8FCBQnly7Dq6JOsHBUa6RP
BLNd274Fzmu8ul3qHXgUXdoiJqQqp7B3lbxVMGdoN1KxzAx9XvKo3QEwkh9606IA
Zw9S1kBs0eiIDQQU0wUIEM47hlQPoGgdL3jicLDu1hZR09knWB0GBzInfacfzBVk
9jcYXOLeKjHUJ8LulTQ+TIeqfAMrur+AO2pXu3lxWWlzUCmiwgB8wZZiLk3jZvNc
YUBP++hqWEp0cVB1R9OKyd2KAMPIN3m2LfBU7r2lpSNHG6NBbkKVf8OF5O3QVKVY
f22Z50MSZpMh6qN+nVNpsyqduvwBZF+vrXah+D0SvtVNra/devZltvO8yZ7bmk0V
fdIpVyESBbWIBk52TVBmSenMa/bP9mcC5rM/2cUWcK2qG3K4t2QrVQv6DRWQgKP6
BeypDjxyL+jqbdjEkH9Cfte7xYPIQZeJyeofbxt/P/cWswH1D+JfQS1Pd4raJhYt
E4fVH4f+o8DvxhsskTGrCXbD/4ZMQsDnbEo/7RY3Pire3bt8CzrPQ9XSulsl9673
XsU2J7ZMpgDOeT6M3dUUOqVcMIqhH7BhITD5cDcxqtcznToIqahh5Vtd1qznuMIr
dD/L4gt1x8PMHpDiO2MrMp8KKjmSK5opjUShk2yXhqgVPr1TN7pnseY1YG0MCYJH
96/L9Gvo53LgiWF6lQ5she05pGngmlLLkSWmzDkhK02qY18oYnzhmFZSSyGE96dU
+cds/h+4U0AF0+ptNFfENktaodvBxkOYa7zEw09ZtHUhsOsE5s6Cdsl/OI6Tvtk5
GePiTizxwOd4OvqTAEwYGveI6JCzpC31RgIGL2onRs5VKBY0b29GC8uzMO5cvcG2
w8HlY2JmH2Ged/Fz2vDj3gbHvshN3mK00zgUJziBYRCwhM9qOb9Cz1UQPx+MoAA2
PZmVEQ6pb6w6aab2ma/fkb3MUxVQ8iLztFyHRw56S06D5D4ATCy0WOaIaY6dJyEt
uzyM+lqc7FwuAWh9lobLQ8LV7i/064UIMmiWSvpQbyvC8M+QnVNcNoj10dAAfehk
AcjVZaZGoCerm+ppgeB6NjssCoNl1lQGst0w5FH9XBdJZV9Enrf1fkrbmSkbw+Bx
/VWfYrLohe2FFGAJhaaPp23BDocg8P/mr5MIP8z18rnCNK8a3pTEv/5dsud8BcLd
0WPIRqU3jlxsTXHs6Kosg7HmBmNJYS3wY3vrZeHuJysE2PotRRf6/yGPp4cvrdpu
1Q94eX50MEM2YBJ/WE56ZSvIVssF08Uq0bnGH9K/LIBLl1toO0lkhDI7w6KDfy/S
lA+ZIh8eeMQq6/UwHWleuCds6XD6o6oHXxSDkXLCPO8RYdkMMapguvsycsIAt07o
MYlbJNt+bfvgQ7EqgWDsyyXg0MtwdpmOam9mDANNc0PxwxhV/e5Z/PO7M17jhARa
+zK7iZ1wk46b8NVzAG54EHmmKXx5JcymxHqGm6Dt3FagPzhOCvCDn+RlUMlH1vBU
1tnNfgZYnokATKxsqwJ70F/AlbfjOky7JGz7Dlnpdn7wS3pjgK4xO/wYdy8c7ruD
vRkSLtWiiUDfSsvDID4H7GBMg2uOfatVJXlaiQUM7rsR1uKSWreYEBAOVvUmq6/7
gQS1FqopuTOokCEr1ewuzA2bwAoV8h1L0zQv0AE3QWNyoIbgEN6MDMpm60BybxpS
pJcTImfmIOiWcbV43qQxrTFXPgTlEDXPUziSeI6mJ2zNyCrDk0OC8Mrd4De9Apy9
CJPZaTCTa3zZ8aN0l09+kkiya2z7Wi69d/2wt6t/2MrH9TktP8sbAHuESNsrq4y/
f1aJUKESm5qWjR+JC1kYFfdVF1kPOl8mQJ2qggKOBJJ5bA0832FNdhkP2gsipUZq
Djph++T73xIp+R2rZNUb298b7wvA2yQucWlkUVvAMi4AU2bLoCRJ6RzSThViK/fv
sh8j1Q9E9ALfwjCBIJrSyDlJHqg0hu2pLk6YWuYwG59XR1pmnoxKV30EiP638IWy
Fl+OR9O1VyzBpadUJC3P3Go0TlIMOvs8/1Dkg0HCUGqWpFAoKwsub/xYi913Wo4g
zMox+IvMESj6t/OtX5TQieizhc+O1Bp+VAi0YqN+F3lcckiaSxKvOWccMBVFk0Pw
B7FgYj5QKqsr9R+IoBRrNMBcnYLhvDwPY2UfIhkkxSOkiCWx1Wt0Kb9h+On8TFuy
WA8z6Xduj+Hy13vw7e6+bOEnP+n9pCHk82ng/uAvs5+Ea67A252Slbt/0IbEQpv5
Tzfx754thoBIQGOE33EVYfpqRCXH+3K7mmv6R2Ich15BhZdGFFxTED00bCED3tMN
zNrgyupjqYG7hmZ+I0v61qJ7qsRsu4bQVLOu5yTpOnsnc1F2Sq+36MCAR+N0j4bq
HFcS2NJD0QQ1YrKtPam0Hxtn+kmGVmPS0r9eXPRQ8c8ifxIfTpI9RtyHMmese+q+
+YmS5H8znnuab4X71ozLDl/qMGp6Z1TSW9FqwcMurKwsy2fbO+Aik4y50Ot/A5vw
iQfO+FrKw1qGIiHMoX6dhsVIEIPoSrxbkb4Lr/jZKfcPMoiuhhTXkVgmYcsEhRDn
QN8RtMhvWNNjzTUvRvqW7wNUplI8Ac7QZKmUwIS+yVicrHS/PYUx/6G3vD9h0mtf
9yHsInonChqmkEkBniuyf6GPBISt13ZVxhtsJVKb/RUQWZHigxMuRo21wmyzDwLJ
zAagQp7OhZAiLuaxMcjrnUc9lkxeK7KjdKXHNMchQkavdD/b4i4+L0bSe+cboxhx
luVaxkRf/UHNQMykGKQWWOIA+oTQkDTmhv55slkI51a7JSkabMtf0aSuntWfpO/X
hEoGAmH2LXLcTLKiHhP7RxrU2JqeMTNBDP0kT4R//GNwiUIg/eiblXyfJLqeW/08
rMi/2vjkPa2tn0G3o8U/LREQQkZZCt0oxu/We+K/dSKaXMAM6PHSJJ2+y7/7Mz6/
CSjiXfOj4rxr0PHG9luaVeGFHT0LDiK5TFXQV/ER0C6OB1z4FWrQ0xdaVU27eZP/
F02qSpABeQa65arP92jyxtiGKAtbZKnL0qs6nTMvp9U5oipeVXNGUN9PSQv9VtNz
I3zC7JH6wLFnQrUvDpvrFDE6N8Txqfz3n3LOHkZUnL3Ht2jXIsrQPHegAiuwbH2W
Wv55eNXO2nfHWdyjck1Iouh63wl9zHMfsRWbfROUGQyCimXyK5uai/aQbnZQT9rG
leplQ//p2YsDY565DgZouCcvU75ioLmF4pI0quP4Ve+o4A5AqNvOrK71gTTLMVEs
Lut4racKYLccercBNifhIvITecrbCCpSvq7xKRp/+0Ek2WhlYafsxMHeLRna6VrC
LPDG/qFpLgO13oYpW3sOHoxIxFHuchh/8L8O2IZzIdZiDKdT5kX8+HeSMuZW6VbQ
vyJ5PRQnZCIMffhTvCaFUEVnQn879LfmrCQV4xKE8DfL0u7Y+U76zDs5nKHkKwXI
hm/MFAuXxWib5gnPzAeWbZ/ZdM+4VQ5nGeWe7ThloNzKn9TcAAJGhf/k2uHioRil
qF4oA8/aBFyPGMkkOvs3v2WLaNR+8JJuHTq8ckK16lj47wSCslluioGc2dbrT1LR
NR8mfHSIa+Yew2SQdkVCe6fO8HCPEHI9iclsE+zXKvtaLVzEH8ccENhlphOTQCt4
XC71Ze911Nf7am4tzmA3mIoB9Yn586OYQKC8LvAhiffQh4fzkjxujvFOgi5Nhejc
R3cslrcThQN+WskLnQhKMMq1VYVjDjLrVCksZt53yC40z78nd2LdPyy1bnyfa8IU
kIuSrHPj/x+dnVbjTTRYc9mHfyadn6pDyTpWuLgsvZloKrs10PNDYMJUPw4DyCpr
gky87icjYwMO1sVN0bIXvsHOYZxGqyD/9RsqkZ53+zaj7G61wcLDE5JgPk/v4qVo
AG0c+TmblfK+YxwQIThiF/JPAqT1aKdoklb3TYgtwSW9OYxkpH5vfYYpRtb4Pk6E
TS0rKZTDMdVMftOGxqEMQASGJbi17P5b7QS27BQaFPxOiBVfYBEJH0q9OXSlb6NS
IsgBrUXSN7B0fpKVLFlIm1jUF7OcIg4h6LeMYiKxTxSdj5PPvzJz8+/yjkLzKEaH
AlZJncoGsjECmoD1M+S8KkWKEl4AOJxNK8jwlgg0ayjqXIQhp6lgp4vzygFIQBR+
x8N7OuOMuQlyneX9vO92hQDSBrotVPZ0kiMrmFd3U7tWsyu+pvxVRjzzxqNw3LYU
hCqR+RKIftTAHPJ+igs9NAm0NiNAUT9jTMF+WoPq7wNgmYCYQrJLsjg+FD+0HCrN
cADh/H9PcdHfvRsl9dsl1z4ZFRoGq214Bmq/AyfDo0fJrsoyIIYQA0zMYkJx8+VH
+iR3rvZLG9xBbbq6dtNJlaEQSCo4dMYaFKbSWHsC5WvqyAuvWreTXemphDVPZGZ1
1AboRfBhzWCOfNpOVUvPuDOgm8R2/5ddal+1gyFKUaVsUZTupEXBRpucABVa2Ic1
rACkNLnpLR5e08j6d2yeCxkkdnPLO/N6oavv/Rp6jqOGQsMxR62LufD8CBJvKUWn
5CrHgvh+Dtq4mXtoX1N8P4lZQ7sZMKK7HpjuENYDOFLcmOanl/w328eDNLVOtlRK
c6NO18QFUIzBXA7o6U3gqATIY17P3BbqvE4pLQOhfCwW/LFbJF39/jlXkj/gelJB
irVUEuev00UYUM/b2xpjgszXlI51OE4X9DOrJdUsDBT1efSxakNxk7LRcqafuN6U
tF7Kgg3Q0I3vbt5VfObLEgrDeLyKgRlxLI0/lzVvZqcVmkjvdhjn5fUWfdV7vy1L
626Di0uMLlyQWoLy12C0HRG8TRM46mw4VZF+Juq8FQkYnO+m5uACcDunSyqALDH8
zN4zlCt9WIqHbG/uOCDAuA+nC5/BE+jH313Ga3oAZf7SWZZwSz5LIwH73+q+PeEX
O1X4nxyR77cH06WtdUl0f5dAwx/PXj1Hz02a4OTZ6QsRPyrfKLtcF514KKCH5FS1
dTHNEYOPzuP2QMRIN2OFo40ytsW5snlIk+czE9kHL9BM3aP/UMW3Bwr4btZSEeq2
60xWcXUp92Yz/KOkb4yvkooaJAILmjZB9vYdkRDnwgKbzHI7YTJrYPbLG9AeFZpG
KTvfIcQySQwr+fHnJifRf6mVrXMXiCeg0djWidng7tZw6mzkc79OdlbE3bV03Z6g
8sDVGsyzJV7J7IkWeYqXkNSBmU2L36KV9CztIsStYt9NnLvxqb3JzOQkTjfGdJx5
oHWBhG7jJ1aBzhtywro0t37JvYXKFTaPv9gsduNJ9en+/rZtf70vcg4ahF/w162Q
vWdj89m7QoTn9d5QSI6LaileRkOczLVxM+i85ZbT2pp7KDbN4ZpKwew7gcQ8R82K
9EjoSwEbcNSKlpNadhjLvoEKz7eHRM2ApVdDb4IvnVT7VvfFr/x0MzvgXHW6pOIb
ziwVphG8CUt9BPEbFnNwj8ZeaI6OgDOtM4ymjyGvSTJtcfxRKN20dzwMX5FzqsM6
5B/3O44Tw1fbtjmInqx+23cVSlOEdMVngk8RAWRseN5Poz7ASIhYcCsUGdGm80VH
Q5hZ8HSgaGwKl1J+RUG2VQ9NZrwOxgFuM8iGP7LVQfw06IbwoaQM7g1SjmN1kUMP
xh+frwk93+dsW3TisnDzHlt7l5jA9dQwqrW2ULqjoEMYUMdn2aNBPVWfbgEM6+eg
furA2KqPJk/Q6/Oig3slQhYNpbAF3Z1g3i9N5cYq2JpK0BUKhXvBoltnMZ75yliN
Vnqa0LmLRzrTKlFseYHnwSvlVv3DNjN5sju7opwRM1o2kLYd35G/OMwLoZ3gT7eX
6NVMOL9m8z49Edla5p6ZHElMYVglG8Kzy0sgbKOFf19t5IwNK4xFCth243/L6mkl
KdOKrm++UCit9iJF81YrXMbCJxwQiYsbTf8gYAliDjpUy0fIOaJaOj5C+h1gF9/k
xHdB73Co2V2TkhwjbiBY0Nu108k+CbXncq49UOSKuE7BJ7i9v6AwTTk0XBC3Te2m
4i4HN0n+WZ1jX1uwWB7uCtLQJ7AzIUMRpM7CgntNXAb5H8rdWeNXygKpvWrTnkX9
F4a2QWrchEGhTbJ/rO/klpA2OtI/MeIu+6RpcdAdZPx3CxfT7fxRc2faDe1OiSAt
Qr65HBCraEVWAsvWdUjx3OHsVLwIBeE6v2istXo75vbjGjfCYPdjzOoPBP2NRz8Q
b8vC5I9kKJv6gu8jeZY2HcUalyecnrBvLZnyAY7u07c2Ec+K2nopD4VuUIzQH1TH
LvWbtIEsxsH19sdek4ZvxURiyNV2n72dToAB0uxTpQ/4ZHJYjtAVPHWsKLr3Aw10
OGbnYMiZGCwarAz6EomPE5REKELQJddAoSVQ/3bG/C/uL7ELQZ8qDzsIpLBcPaZ4
2jaet430FKHB8VRexzxhjm1tGdjT/lzsOcp87pvmIoq8nJIR6cgfqdOhlXVQCv8c
f1ZU4cfz2CN2Te4Jkxlytt665Zr9m0MvqrjzDQRJF+rd6ZN9IHOoxXRcjnuuGj6G
8oqhj0IpNJ+bFqjO5Tt3XhgLSX8wPsz/giCSFrLIULEP//Y6RBJFrXfHv8Ytc7qH
LknGqh59KpD/aSGrR0vrxhz7A0z+0jI/DI+AkwrMP5dIatsxnisGN62hvIMxa2DS
S84l270bSYf8JLy+uJrpe31SDziXhPjN0j1/z1gICs2gmjDQmSKflJgdNTJh7tPC
9BbfhTGb9KrDiwC8zSKPffaRmN7e6zrW6Q/7fSlIApc+ZKRtc/0B7Xqrgkma2QH/
KTCa1U/MPytvW4b4WtOfoLdD54WgMVO+Nd/GRgkTRQAEAtGUh+gT/hqaNp7XzFpS
UgNRicfhFObpFFK8vYBnj5rigwa2FDd5XfbSSHiZRUQAY4qcSXR/G6ERpM/WV4zV
TKJbk32PSOrnGbZZdpqZ4BNnOtlQ67amTVEeca2vX43KzvZ62NEJ/17t+fTF9pC8
VlSLreGf5WktR9BLb4GUu13/E/9xSjl4VOmV/RTY9jgwSgXSZJnLtAFJDWw64VDG
PZysKjoJ7LIUr6IokURJNMZlDR5BM+O503AvhJqw8YXMw1YQMGiIj3SP2rmScDSn
kaYCbOik1hciTNcZyyzhgXJWBD1831NLweywrItkGJWy+CodmJIBnK4vQYQo9Jlt
S5u/ySpv7IB/6WOdOMNgOPWGuP4WLKY0ou828mmWVonGyHTPX6XpDJdCCe2uE419
Wp9C9FUSFon5Dxr/iidpE/oq9iJSI8CCL6dBneSghmqb0+t9whqFykCPNsqr6SF3
tPtX+BvLs5TY6KXruRGgODJS2YJjPZnDbAuJ3MuSYpyA4ELXQyNUpL4kLkWWqGMa
ztPUWUm9CC3oawR2n6aaRjx1m3IGocfqUzeZqMPEnPFCDXB66nGHSb1hUfhdAXgC
dDRK/x/VRLdejxq7+cUyRw9sN+PMWZw7Ec22cnfbQdK/EDyYlO+KCG5FUouNQg2S
h0U3Uz9qrsKciNTiS2q0OKpvFW1Jo0R64fVxT5jw3jyxQK/YwyNLvTwnFneR09re
g+fNq/UCGj/qJhRWPe4YD1+ehAVDDjVUE52VRQfW64PeIkvoZS/jtabkyo24X7J1
icrPadNw8VT2kzQqkPe8mr//fzC3ezC8N1b5KnWJLem5sD3LH3hiJV45xi5ItjD/
eKxvWoEMau/sexpwt1uys0MbQmie1/0dqF2hUQ9CX6HaUMxS0eE9N79HZRzsWg0q
MgHevw2cpV9KZcPNXDdPd7rMcu1Zf7TPBxdYMHLmeBHP4KTP14rIoPaeu83QUtoX
Ku7Uczk7ptgwvDjNYYfL2y4hnwSEmp6uvFlMIJv+IqDDPTkriE7r8wkotMsX6ulc
l3jgNCMZyp1KXqCZArifgvAh1lSBY3BVSga1cURYtSOlkOH1/x83ITG408TRsDtb
B920odY5YSWNBD27sDsJF1L0hD/yxeAfmijr4BV3vCVXpcSmcbz5Y/QRuNz+v8vZ
sJumtTfZDSsw+tdjCV0lBWVYvlQEuy+Km4aBhOy5CWIClMzEd1Do/PoymZJLuZwX
5t0vHa0w3Aut6KKS05ypOtyBo+4z+dHc8boQ0iQG5/EWZjjmu3eDiTqowb73wsZZ
JzpnAxGikqzLkvk2OAME9dfP1OQ5cZOiM2r8Rrhb3wDEAv/AgKSA3BKHiqNA9dw/
u3eOo+pL3BnFOt7+hSiaJ+f06XPnKEO2U/l4ZghaE5ecZ/WVTeHFIHgFVHIh2EBG
tfkQhhSappNOajzCzpPrzGuHBLpNi01EYjV5X77DK6ZghAeIXlo2mwQCc1E1vStq
huznin3i813iHY3IHMVXAjyhXcZ1TG3/4qYwMd3UppcRGuFfruCscIw4JydGCgj6
3DDCzHItHfM1T7nPV9DuDHFgnF4/BTGocqBoDkhM0wtj0HMft02nFAICIMeBJGW9
3pFBBVdxkPDkGcgyRl1bK6ZnK9uRwyA9Fj7NhvY+Dw2jXZg1zt1Q0tFxbx0NblTA
UcIQ+M+47yxUPoS3Np0ee79ykgGc7mMXtbHUOLE6iJJQAXPzNwJFv1nqCAOgJYic
N//PHv77lqfU+OvlicDHreNdq7A2eC37O8xmxUT9gNbfZ6wqFgp23o0QQ03doMXO
WmgYlJDCxkE3RbziNXodjjHXiyT0LkP6kvZn6pyqUwDTN2o6eRQSHYTTFtKc0Ndo
84EwCaFFAu7YSH/wc6Ongshugy5ASXtUdH1L26SCAKzVBl4sYHI+Y/7FestirO4o
IE1LoAPKjeX7v5Tp1SPFZgx1w8yYF/4LKFDc2p0JS1uq0aDJqQddf4hvCru/rfFs
spvLnaX1eGOUiFA9yFoe9ENELuhFPRUQ4v2rgVT3DUjKYrxTEc/CVtcTQyAGkPfc
PPaAXwAbd7C2+3McwzPeg9g4Z/ExXm8dSV2Xn4C+Gwu9lFDOEwz380+IUdHV0S9M
gdTP4m6J+9UACFHPsg6TPXq9ul6L8rVngpKtoCK3TbbWj0Sbw5KF/X5JILNQ+x2l
vimAUEJADD0+Low9mao9e+ZO1Knq0no8fpPm03bhnmZmrAfmfIytKHh6f2D7pwRG
eYA3YBo7PzErQY/ayW20jf+8nyEVafqxnCIlCH7jf+Q8FNlmi+NoUM7uBe+J1amh
25wQJ/v0nyQatHUQm7GFNNv69OUrxO7jYBMQT+qqGO9OXpqjurVh9ciMRAfcg7No
ZgUHZ8i7jgqr+eGOudDkz70O/mh4GoAVJNQ3FLVJz/owlhL4pTDnShuyXhJqO2Gu
41acJY0qZZLOSJAv8nWleUvWDSfgBCguOzagLtI1WUr8dIwy8iYnOIc2wX4h++ZO
FeuR6PA5Ux/O1brMlAPJk4T+apSshTTO7a3GTuS7V5eOTwax6PXJU3w/VakWLzOB
CNSxl3Jtv4xKeo5PYEahZIhHiPkBE+7GDpTr1vJS2b7neKAsUuVtijC2xj5yYOli
9xo6Ry52uoBSTfPI60F59BLxM/X/i1a9grjY4UDvGfJPj01Qvo/IY8172MZtob3l
NaQMbnH+tLqq+BNb2e1U5ywzFu7B4LN57KK09Uy8FycOfp+Q2HMjPg6jY+y2x0Qy
xHXw6e8wEbHODL6x3kDxbnHCM3aFQORPCqxeU4Rt8I0fhzV8NOHjxxQf5BkC7eV+
By18W1LQ94om+ElSRgN9C9AbNmVQt3in+eU7BXQ+PwiSZvpDpZkslkQLc1+DOfO9
v5x2UX6/FS+4WWSr1fjNucYmd5Wx/IJIfdfL3YqrpKkUrXStv1p+hfN8URwosh5j
q25TblCO6GE/rugZLCzvehIaQr45+TQPMTMFy7Ky+/RuOQbaG2VTvRSe0aRwTaiV
j6gtF+LEVYfxg87G7aFbN3lAmR1KtMikl9vs56K4AHep1BWaeTW7zdM7xPBoSTnU
gacZwgcTBRi8ALAEpX3Qj9foR7zogkZFGvDOIbHquMOYDuXUSF+v7LsRYysRBzRn
pJeqDPagU11eewvZ2eqLjUYu3mTF9eYkPRnJnnveekqUV/TuqysvCnB3sjA4vBXK
Fz8s+afOajmLQTyORLNwMuOU4o83YnNPNIQ5j0IAksF/WkPlKWzN9w1AWYUdQ9JH
G7oUiGUaY+3Rt6JOE7YPZ3EpPEs8Wgdo7QVxSf0JLYj68E3WWAzGnQyVlTsptMb3
z+2wpY0LsYlwFDiyZPTSpYF9/jVNRawOwWCoR6P0XeQxS4VBiHkWeC9dh01T4Qni
5Lccg7QpIhv5d0x8sVpK1BIveGif4Ys09CJ6wH82OWBme8X0QGAs7v5qHnZ/Uesg
xobEill/L2vnfEb6qxXWA0ed3/gloZ8WLRpL+xWpbeQtjysXuifAGJRhCaYWrvRO
zC+xrgXSDWYD1eZUcWUlsO6HfWcn9RZsHDs9RbbxkPRa8TkRTRVZABKPv9H5rca4
+rqfvBayJmMFoWB9OKEm7SaxdLR2Rocjrf9bIx8COKlwG992YPafCqWdVHswricS
rPAQslP1df+L1/lddUMXKJvdJssEl/HOb27yWEs6HbKNZV8HqoYWXn1mT4Kafry1
IkPA6qOnF0nGqs22pdmsUbGoSdA+uE5y4+jGFLXXCxWGg4LWXwQELtikPjjCaG/J
7l1xtKqkOxluY0FpX5pPeqAdKwmDdNvpMKDo9zR7TgBCaJCRuwarCUl1ELbv34nW
ttybgCZvaXgJbnElQgKwJTaTGzoWDfHfZisjXJ4lp9vl0w/9zFNHcVVezFSmtG6M
kMqEujkEhtAN3m7ClllA/wTx+b/Uf50FRmtbjxIIDADIgbcIgmXrRdcP++VO/tTq
N0ONcyhYfN9jArG4yDEr2XbslzTUTNNZQq4j0mLkO5kCghlJleaIBfr7rON5gS8K
t8IcDRbVCpuT1WLnBPiCIKBPgH3PNVW2xZnlQk47je7wptMHnrysK+rhR29GziI2
ABEuYYdORRJP3Tnuv0vsQokbQ3wTNDAdMQloy9erecxFEjd/3BYYQjxrlF7tbqfq
MeA8HXS293lvSFeKM9IEsYkFaFttfTtqH/qT9L85gIZjdvoVPoF1CO/7aRxnWpyB
I3De3ssZ66P9uJXRk5JV7/pOIgswF1YYQyEuYS/+VW1CYtLep0HSoW6814D3n+cf
/zp4EzAVB9qpMg+6HBK7uA0hmEo65CXTFiyU6PmOFqTO0i9llm5Hhlu58+GFOxbP
vmc3HrvlnJrnjFfywguxWewt7vEkzdVQYr0PvDUjcesTOgmo385uGv7lMPXnexer
ZZtlQNtdCZiPW0/xpUfDMjj6on/WVDaO9RkGGiverjHkTrDnd2JW+hZawnRxmpG5
T9EAlnpNHdLML0wpO++s2d94hFU8RC4IYb3L5c6NaOt4nROwfTcIVKcVS3IT00hM
68vHMfKcuVXKQW+DrUo1lMpnve/2F9m5ZMV+XdnoKSh79r5GWPP2Xt4hYgHvs5bg
SkfGynSMfBrXtMy2kJohu3vJ2sB7r0mJcivU1PcDpGDXDbZRS55txKdqfq7EbC19
XJjcqsKatGSXZlcsrEVmzXEsVVjv15BuGzm2oUXJGND34jAQ54MjXsTwgCXVKUuO
5PC1ZMhJuUVlwQBHB2TypacHKqxY3GtCYUITB8wGmbychTeOoYxPZbLxeIv4d+X+
85TwL0b+Pwxpj8boloEU3DiisK5rnRZbB24D2VH95q+ko0qRD/xSZ7pA10xNs8GM
QC2FSpo+wKxeKkcLLup+JVrEnPWlHyPfaXDmzGnBf8RIQh2G2LkKHnI6ZGasrLp3
14GkAXQ/XX+ZcykyeKAybVk8SQX/TBUHHmrC5FQQ2SEopdRRooaznGaslb9wnoVY
eYcc5eco3bKowVPX3Ywoqf8QoAUahXqpPIASW5xuZhy59CY2ymvSuXGhuRkc+e7r
46NRjdHRaojGuyXWWxViPj+L333ztX/lX+0N2k9A67LBvM0fkunuBIjKu67Ye/4U
s+ZNC9QfMYxkmhxsrnM43PM0XLPZdJ1yCQbQRJxx5QSJKRh0HbVn2kYGvOrfn/DC
9NHbN0hHs6X46KW/ajX6RaMVmp1PDQCi8PSKUuhiEcwnGf1QocMVSWajuZ2BX8lB
CmsKs5beKxsuQFLq7OwGX3MRgmiAOhpQhVI3Txx85JNZAp0tikfi6TeyA2Oh//eS
gYsC3hfeLykVMaXpsLBK+l7ZBjAod7FZJZvffffAKuW2c3/TTKpwDrw3RoRoh58p
dOmExHcXjYnk0OGRC8BtDV1rT438wzvytt9/Ob/ELsle4vQJPchndo6DZ1wcgKKQ
w4K0oiXMR6BeqahOUexahw7KtFd+9k1CVMgP7Lr6tLdE/1BGoQByTJq3Bl3fDuB6
gE7jFAYHvw+MHlmf37m/hWI7ChFXzIKLhSvj+SyveN81Goudi2dHlFY+8LYQpBPg
C20e1KVCZmuAVv/joMvBYoJx5Vw13cBbKwb8QMb1LCxretvT7RDagBY4jttnhWsb
wOFr9Dx54qy9BrH0G4DdRLVde1oxUgsy7gKg0Kb1iufZNEOj27wx6PIIWqKfOHjp
gEz7a6svT75LWdXdkY+CsRdcyBGAV53dwl6yTPqHQM/Cosl29Q1AaNS2QhutSoDr
vZC+VQlIn5X4Ji6LpVSGAhjfRsQsim3eIFlNZxvkMFmQ7CsHnsDMhFs4jXQkwoz1
EITLKz3vGclJn8c0T5KGirF2yKBV8RDWRMgf3Q2jr7OPX1AQhC+ke7t8gyw7BAwW
RKdodNB7AhZrPeWb+dg4O+/UdVTIZWaJymqg8m2hi3zTR2+LOlgxWtOwEwgCtdKh
LWiOFaMWCBu8QMj1C/dciugIwc41Yck0il9jbmj+990uBpU0pb9n/zsOUpToDVA+
vJAjMth6lTBPGh+Erwy0wdxbg+EoeOH32O2nMQz6ko/z/0t21q6UsJPaLnkYailG
yyUR5WIl0OnqnGDSFDh4FK7XbPodfyweNUUX1KZ7tb1qUBIPSMkhBonKOxQVL9gd
iS8M7Rd2e2qha4QYsXR8AWcTRzkSzXlIxLmWS4emq2zszLNLBCIN6d1WKzO22At6
4dKuUuoX6+0Ss4+8bXZvtyFInMOpz4qKBd/vTcYWaToNmvEzpJoKOEf0BhmbI2RG
mZ6trNnhfmvx7iPXBPFKE5yEtgrlr4DSpakrcwtWbraFgRHyy9DkbIizLeXT9E9o
27VG6J+fhjW25AGu9rwjDuKEqS7TohD/pGrY0e+4za6iMzZSR9hEflwRSJ96texE
xGVW9sVcMXwAYYCEdB9s8zvhl2N8HYD/icO7KRB0RriU0EUK2dibfk5cWu4GlXp6
qLazK58edINP5sGMU83xxBOvtR5so9bYgfWvmGD02ou+KJidBKBJLkBwabPurb4T
3G7cQGQuWHLevV2zrP8FNUXPJqIjpHFmzQ07jYD2VMcHIgxhc+8hhc24KJUs5YS1
L5Vmp041mzbkX7gJ3Jh0WiuwGty9K/MPqTDJ3ogEQq1bg4vpPbycVtijsSFjmjYg
6T6ktchjhjEd2r60WOBzBhZzIBO2y7CA/syqOGppkKAUgUwRFXuRj1LBfxYbBPyU
UnXK2qvdewxtVUEAcJGxfokLAIQUweqB4xB/2DHDJLPUQSzHaPPtDA2uDy+gfwnm
IgyKq5MrTuWqLTCtW+iGtdF9t4WTY3DDxtgkjnQNvwI0Qb6kBNX6Xkj/muuWw2kL
o6Yof7DhdtHVYg/kdGhTP0xPAhAtdYfVKSbF2QKkW2/aI3QAe7Jnh7J/8/4tp6VD
NMYcELvlLezEyApskiIbdPFyhos0vAMIxpXHFmS81zPN9lUZ4Ywf/BjVyq5aJj4i
/Jk3Q0ve1WZ+LxZ3pmBQ5tf22QR95r1CR+mhUJ6tpouqnGMGI340izOADguZZiYg
LNBFasU0BfCrj3hPjJdO+j/tnrY68jbUglilfNIRPeVSMJTGNTZEQCHhBxOqw3mF
e3qxmVYyPcLNYwKT9BRyDdgsCE02m/WpIOTajsPj/42aVRrh9iae2kuCWZgN1Wez
Oam9+sI4NzlNEpZOEJageEBYSPkt3gqWWK2CelQXws8UTPjW4+X9fR6f/R/k27nv
ziLOCW0dQfyY7ot/dNFlY9QibJaQEfLApzBz4nVCBWfdfvmErn/Y3/IRAlUERbeI
fxUIi8YE4KO4ILiUckIjow5kioGAhmsxBh87pKSuGERa/2j7LflXiJopo539RuJx
eOYBGWZN/4nJgB5Yy7nVjvtplQIwBA1m/GQU0oavJlJ3o34FiMlHIQFOiUD8a0gm
MoI6qAs5RmEN/HOT5oZM93PY+QaWVsRuT71dwfcFadMINES5A82Lwbo63qq45ArR
rntLe94x3iLIsY+AoKWvziY30fk6XyHt5j8xuYZ1NmsVl7FSm1dNTnACATp8hf4v
71i7VLKqns/tMDLXUO1Kq5xdcUVq30HlC8EV8iF2sQ9RRr3AVkCkNxej7JGkaDKy
3iZvTd8M4bska3Na++8J4UoBJOjqmaxWEuUWPj23uQuoZeHiNctmCZP4vs5xFS1K
PNdGZ27oT9M7QhkCYw7tIT/csy/PLW+nKCJhEstHt5jdVaj44t+a2LNA6FINJltV
uM+9IhHPwVMbznhRkYYZSBYBnnuXboUAatsslnKtMLBiQzs8IKrhlKijE+HpdtQ5
WsG0/mq7Q4s9HCJXBM60NneFlyjeqPya0R5D/K5orGpCX5BrIB4NBBYtFFp/3lS7
th93HwCOfdQsoOlu4BGAGcDDwBIPbMzTVOzSaokXlcTm/EPaR6pRg4smNsWMDgiz
LkF5DCk9t4atAvXEJzGMLi9IwF7ejKdRVW1nA8xObNM1SQ3oA9NXtEcG9cHjNvJV
qJc7OXwCUGxL3sphnkVUZ5/Edq7+uIc8eqvGEEle1b2ehRJvBJlzfq/S1836xn8W
R+DRmzkyEaLvJhuXsNdjxUVv6eYlUw/5XQhGyOA2rWh+QPBKTzcClNdvlHqsjIPk
HwqsyKKqen/qkU1Dk5hHkgcjUHgNsl7RzwqsD9F+KybLAxQNb5sD2hSHdjkx9fcw
OpGaqQ20uhQ6WjOQGZfW611X09rniMcDooT+IgwYltohu9kuhbb6rc2aDB2RhPWO
nQ3y4vlBsuZ42yGUHiHwH+1fCMUx1Y2iR955N+Sh/iN2/UN+4FFY6ovZhIamuB9h
Xt5yTsLzGbYgrKdg2ysojbMWvIKyMmqSIRaklBnDSGHzW95Og/fWN/DTY+NbiGUU
Xg6o1Ebm5iUvLvjMLpo+5PgPtm3rs7KK1+hFYgmbTwJBIX0IYvoYmCS0AInHBt3M
qT/+ULP3AiwNjdum6OXfkaXWQK5PVjwQrrUAQgiZrlP5SWhEIAjLnJ5yf6R8rcCN
8PLg2o+Qes2G9+YdyeAKvsD4N1xGxIKYbqJ4bWr+QDXl58VLl3jmEX6+No7YxtQe
jLqRK/KPNiUStOUWCmQUndFu9QaJ9YExDELKgsQ7ApdsufznRTGRL7RBXiO7VaWO
Pw5ASKrG0U/BHTM2wBUgCXVIP1YKGozVtkuvvs422pBIgpRuWz+WxzKGZ1Mm8PGn
u6hvgFaUINo09TNdJqpd/JGb6i1hA26zltxhVIZMQ9w8o4hTxBx6Os3SanttnwiE
bK0cPS/ErFaGY9lrx7nLfAJVM4qAKSibZcrZrEGBlNr8KLj1mDqB9muCdrzpLwLb
HhYbX+cyej3tTvXTZl3WYaqusxaXHwHti2yChtyeXmb0ZMRMYNhmvFuy0kX3FpTY
OR/H93XuHWsJSBPzyuyOJ3Mg8nJbeOG1+f0ELp84rSDrAUyBCdHQpjYvX+vbjcgC
826ZnkpfUI9xKhS/trA07kVv0kdS7a1r6fk9cpIClkZwlkzn+V18gv/nJWn/0aHJ
IcuxF0ovzGF0VPSL/M1i+HOYoU+Yq40Qsm8hGZYYa1UryYPZQ2YMVsQigWH8uxEj
xp5JV9+lnoNtUC7kgxfn628i7OomJMIqYNhdzJmXfLaHFepxkH5iwLqtoDj/xYiV
4FT/wlg32zqIL0ZZdJFJvwQok/92Wc5iZ/KTHCG+ANEyK55uOgS1ePM9e50eazeq
HlV6bHN/y6SYDrr6fwWYOF7vFQhxkRv/z5G+EgmYCJhc+0Gq0gppfXLrv1TnTv+b
qYwqbJ5GEZfVKdQsi50GydcRkeg4bLUQDIrPzmdUhnvVS/z9h5XYcykgPcuPvwuZ
hzYTrGilGJbiTrTLHp0xdKdkvbXPdAHIiL9NXHUdS6zOrZQCe0dw0CIvUlIyE94E
UqBzH9cCnsUhIthdV1DgiIkFsVMw0j0HH+zU059EmJY/Gy2/HQYCMjt82XdCh1fV
hYMSen4IiUCwzYIS83rME2kUwHYAa5I55ooQTFypOi3/kgVWE7It0JgATMW7MNX+
2lUvVs2ISW3yKoNgsOUhI2d4/rWp4vv/qhdrsVKFS92Dig1ehS0W+Xe6HZWT/OL9
+UG9dWz71ZmpRppzG06jIjaedzyyGe3GPsc04rSYT7+eggL4R0cZmxAP+FwNaN8n
nnZLIVguk7BVF9h8o25QKzFfR2byb0sxEzUdPLwYt2CGvPBi/ToLn+Ar80yhHDc9
IrrkqacaUl02BmakcDxU55JkOy630vkaJdpOWcaEFI26d/KRUQDaCrxsElG93/pf
rLMdW/QphwZLIBWKkGD/ucPlFxrc7KZ6Ea8HvaOHEFzlDBlMerblLD+agqEKHUqi
5bYc5Ri5E2ct3kc0WqylHZ3KJG/J7+Y/gtcPFQ42RhjUHo/hq7S53IhiKt6HdWgF
D37jJd+Hl1TCAaKUfGvrFwa/ikDHgh3+IhGWgR0ZnwkR2OLQcOPsCsqht6l9pJrt
mPtx6BlIKA9heq8ov8STeEYR1I8N0N+oywE8QzUc5fYKE1elWySqEDpD2/6/hl4i
Pv3qSo+oHM6FUKw1Z42pTwaq/74e6iIVTG4WRksATo3LNt7EDMBfkcoRUFxT437s
moX+y71V4qoxaAnC9ikuGKM6gFm/jHEunUdOmsU9BlFAuCISiwbWHrfWwlMEuInr
fgE7t5u5IxeF7X0xxQ09hwBUC9S2R98qE5HkjVBDrasHYINDKeNBDXqM9Lt+gfGm
NOMAbvYZ6MbIcD4L+1fH1Mbgc5dtTOgue8BBBf5W4JaCdBI3K3OaYlFogyq1fuen
WyqHchpGC+9DcwFgTIpVoP3urpX2VjwVrnOf+bwUFJ7XVsG47WmIbHxAlr/6JMrM
/wWd+8mCliLDCooN1DM8H7IR7yKbeR3fLGdqVyM++h1yHCA5/8Ei6f3JtDUv7fJ9
dTDf35T52HWMoPBTbMwlt6cOx+UWd0+iyNjrziggpuWaR8B01YVi7a2UkFon871u
/G2nOUPYWZIdC2FY0Ke0cWb6DeEMJ5tAAWMqaGQaHJT0foqGEWbUtokcFQbLRWpW
2AY+qmJIBL8+wHTgUtNtpDh8CLnQsyncpmroFq95LrlAtxRzs3jgKlYm9j3t/zqb
1k40BiD3P9/kw9HJ1GVb1Y0la+d91lZ34nA75iyl0DBZilLD3jFNPth+MMwVYXZ3
Rf9dt1mD/zITqX+lvknYS0a0oORDx/0x0qVxBx4KQQ/w6uXlbGMEu37FgzoSvt+T
7MyCCc76ggHGOrTgkolMOeCunf62q46pyVzX4Ni9A566CX8FJ3w4sJ5nUBHD8m7R
I+oAD4Yz85SyuKTNxUb8DpxW5hPGFsx35NwoLpN/hhpWAWvgSnj9IYeTEEGWENYB
3OjQudh/CcvB6nmn/iiwCqALtWPYu8QoCSKvd4WHEC1iUi4MDtj5qT+9Spft3YzV
EAhox3siDfciX8zCPY3THJLpKaCSyqEZEchokF4+NZ37YZ3a0boUwoMWnqWDIfX0
p36z3ygmkVrFCr+XxNsMInAXw4wBhQIqxAPTktUutwD/28uXEJzP5ccOv4XB/jyb
VQNxUSX/+kyVa8yay+5Quap9byGRNH+uL0XWyb+7D+lnmSUEmy5+DU1SDDVN9Thr
ngCPNsVb1IQ/S6pxDXCtX5oUoIh3zluxQdBRrJlYWa6ak4Y7dQ/UR36njvAPZpCo
qgQ9I/uvycWaFzQcNuZL3hGS2gNwTLXNjQtQ8t0ZkGIINejjPIAbka6yt7aBP4bX
zlJ2XhjyrkjYEeGmtQBRjNSotd3LHTnx68YPI+TTT6fdBYawZVf3HaU71Rrgmd4K
Uo8zPLBNhDV/mKpChqrh7Tz0oHOg/qj9IvCnjpMHg6DKctHdsaQZPuBPKzlhU5vP
3N9wdoFo37nSmvvPgpmldvG3HFEYr0JH5i/fMYuddH+ntrP1cJga/CiJ/9q/RmeI
h+aoJzjnAjiDDEcBW4GosJ0Wj1tXarsFmKa2llHDcYUWN4XNq97nuF3V55gzyuQ1
Fvh/mDWDjcrilpcFpyBD2TdAPXAZdx2QXmXo7zH7t2ZDzSzhb8pdeTIsKF0Cjqen
2LhaRyRdjHcQ/XSOhumc9P22J6VgOGek3rLZ7lfYRiuf+AkJ86QR9gZUUTeWYHrc
qmhSX0x2moA4IYRnmdHw4IFC5RaWSp6CWp2hos5Bm0OAC6iZLtjaZvsXNd6Me/AU
bWpKFlxuL9qVdczk3HQ7/7GehXQTVT8RtdSjQikgbS0wnATev1EsCzg8anXrey2S
3ezm61+2C0nP1p7iTRBFDt1OcM2pX4Vwd68vlH2KOAzlL5EvisRlBxLpIHShrOC2
fufNfa8mC68q+7xk81cpXqddirur1ZSs7XZ4xejJM29+Bee2Q64tdF9Q2Ko6uea0
vf0S4OBNSL1xAAGtnEkzJ9y1dWOXGxNN8nQDls4DNekIc2hGn82d2jcbisaBEdcL
NA/v14Lke9v1hQYlwiLV2mOzjQ1ccvgFmVQzdLUZ/v3nPypBbpdvrN0XkZrRHOox
Vr63b77IHoScNNFBNWh9J3uA9soBNbBNqwHoTt465zDyJH6lT+rU6h/45FUFQsrN
9KHoKEyeUi/nVdceFHwOJaxWR6Y9lgCyBDkP5Q7aAbbWX5jscT7OHgsD/kGZ6LU3
ZBtNulm2KnqBT+Daju124VuvubqbzemfwkzI+YNBA7hfl3CG7ra2L+Yciys5kyhs
O1ahXCmHgRMaU0cePjkbtwtn3sXZ/Gq3EKGbGnMYYmpS+1COF1xxt8J9vXlxilYB
yli0YfVRFzATdy4vWj6uNupQo5r8YaRZS4Kql8IPeSIHI/U3d67p2b00vCqRIzD+
nh3KXfrd6yXmfORY7MFYN/Wl/UbeY5XVSSB6BDrWD7vBJHqkoUE8n2+DdPCvZKN3
rY97X5TZNlDQSMZ83onOpAOleAvQJuJiPDrI8VGR78fpVHDdSc3UNQ6xhpQTu2A6
McqEFNwZuXbz99aImxb0dUIZ/sTG7jI/GSSaajxA/mFu8jcGeoRd4SIUl4DQ7YJy
r+bL4hBIED6qMCs9mqQkLO3x9XaMJJH52olZo8gvaMVuMEX+Jc8YKeJLf1jFkOht
QhIIVUfvbXK5x2clIicho+GZXFox1yjBWMVEYO4f7BMNso6rqIgjIMesiSSoSIsz
b4siraH89iYxV68T531/cS136U0wrsLgHgWHH9F9GyGh5o5T6aQPKfvXx76yFMJV
XHmOYfBeg+VAAf1cl8OIM2P4xikuldqHTrlCX37vKByU1YHlhyKkD2jePJhGcTSG
B4k0WR26xrkPt4sRBzpnEVvsTyiUeGUp0oQS53pOFa9pGddioVS/v0nIcZKOZLTq
AruvvYCWTln+IY9Hw64jaezYIMfeUSUsCvARDPgJOEC8H7aLVS8jaYSbMhnFwTt+
ojD2DmNy9QZN8NDA7Qq34WfMHR2UtAqahuftrM2rE1El2ltYpU1bbuKgoyRv1Ukg
sPMXMd8pzmtOau9q9oFS20akKliOBAHa2FQSPOM+MqFE4FFnVd/fk9ekLwJ/4cIE
XR2iU/GcKfT2zdDxBGzU4mMGX8pA8Pjr7Ce0ghhzD2TgdQ2M1tjB4FgCPhsVt2a/
yGfPSABZ9OmDBhJpWbGfa0zO3gaobWIwJWWLwIiBisRysm8Nze1F5NV3fgREk7k7
YGm2E2T6x8FjOu+thjRWxpsgDfcat4AoPAbneyytlaSQeRgqR82lhlVChdjNQX4T
GmljyKni7L9HIMU7lhYrtr3K28RdpQMv91Mx1oTMFDg2bXDzetxfnCPb49AFZ5+n
oi8tFicTWWd/6YrVBL39AWVKHAywOTOpMmkzilTNPpwYA/JRRnb9+Bdv+AKrCW/s
MEde1CDdW6a5wNrisNMryPz0fmNKtWstbXGOq1Bsxoo7BUniItOws6UKI+yKe7hN
9nZd9f9QOTxjmQQuHtI7PHbksNVKJJsZpRXVR8n9pEs/qGyC7QEwDAhIhSj4FLkx
qmswO2zJPj8T62XW7yxwtkestHjA7H0HHpdQjtxNQPYFFm4+fidQGks78mmVTEUX
9j3RNzwmAaHMTvxqCPYwEsd7aVvCrKVpIWjj0kjJKaT9COXVdPVIsp9ZxYvpfQ3f
YkZdV8mjzMraDbzVidcapAvZd49bhORkJUqHX2HmSa8Vxu1CheRQKdG35vTBoyFO
8TdZO9AJQ+R2SoUmN1xNon+zjjjjVOY6PFz1+xK5fhjXGW32TnvDi4aTeGMhoSu3
uPHKzK51PYRsAe8IDAfnaZNzG98wWZZeMKT+dEFfO1v1zunkoJaCjGFzTamzt7kJ
vIU8TM4CBzJlVnySaHTXEsQLQDFd+3WvJdxl/mc78udAcUz4SPav0f1/Qxs9pfzC
Y8hEXFMuAtow4wEaubBM1n/HvI6lozR9Maa18HgtpJGYsTB7NF1W3Ar2ogT/X2Q7
GwpXDNay7ng+bSoGc1INiS9g3wa0xaNi+8t8M/Cpx+Jw5p+GaXQaOga2MuxxkGTH
FvlmEwFU9Tnj9MuHqRLcXWNAapsEdgSTJBHvNXZo+L8/xVOBaiHfqMWnzBx0nT7P
XmCxmVA1Vbd70YRKxjfsu88IglQM8q2M6SMHzgtcLX1ogWn6PkInNouUcAZ/JYEy
Dbq63TBrJbZixs11nSfhCG4f0gD1dDvQM9w2aE4YeX8pnIgQqkzkY5/OPU8+9zY3
7eOiZfRFumpSSf74+siYR/c+kRKPWpvXVea2VaOTAd/dU+9GWRkA64gxGOYDd7Xz
y72WUka7yQ91oFSmzYB/eP1M1mkKUCXgOhEmF4R2GZ2fdr2H+0+uQ+FohzKzUzAD
HDgW6/+VvNc6bIqtK8vg1MWYQ5+sXWuG22tEcVt3hPbrT28rIndYjG4jMFfZiJz7
iUlSDEpt2xHNvETNroxZ+zwYXxpxcuwK8tigkQ6p8rE/w/tavBiJBXmZ8b9+nNN2
9+C5FbMseyrWNAdH6JXdkfcX9Mty3tVUdDtu4aGUWpqQ0HnrZ0TPG0AehMIzYFOs
JbLzNmnrj34ewxQqe5Qo/O28y6ld+InHqqNec5ySizKEPYQ7KUn3OUpASHrSMTvw
SzIHtb9ucSJiU6PV7rs8xdqh+nPL3bMVg6bRLdjEvlkljDGG6yqHQl/GbStMmX7R
JWHeTTz7FEcAPXaG4uz9kMKrfVy09wLieeGkWc7RCkaU/dXsutaYwAz6kZnoR9uW
jv6czcE0gIJ+lSJW5OU7wCmghL124hZdjPjfIxA8UVVee2e5kNy1rhf+XRDOIBpw
6MIBraFfeg88lnFUh3GKw8xzEPY2Pw58XLB7EqHME4bblDfMnAM1Jma4c/L9hHxD
5TUMzYhaR6BtvKzT8aD3n6PX1mFCFUO57LP6OOL42slbL8M/Yrhc0nYl3zi8tfuI
7FjGcy1v08qVKklHmf+jkLx9R/6T3GCfYfjVV3bdJSnyBU33wFRh4viciUshrXmH
vgDAlvx/0p3HsP6UkMjk+V/CJ//uHEqhp8OEXgy8ZHsU84dp7EJulzWrTfsKI22g
TK8Q+pC3oI1LkSUvLTcyb4fKAAUpZRWJvMzv5ah50qnf52QlIovXEBZGTNcm9oQL
MdaEE+QsU41TIpI3x9uNd792yimwsX1RXF7WrA1QNd8vrxD/DChD0paZgJVwy9Ed
mdDOtPMGgdKaY1I3T+mSNQX4gI4UM3Dh1rROcnkcnc8DDrldDYxUsSiMuaPazmV2
zEvZ/000bQzNMxtHM3WzdEt5Bpf0xrBQ8tFJGQWz1F6dUBNoXl7Nypj3D0Q//e6b
ABsG250lKVgJMHks7B1uC1GKhqOYl5N8iablyiC8WxEgu4W7YtHZp6MxHxUjz/52
xtuPwSwTfEu3MKiVG1L7oVkLp89IPJUEMxz8FDVf8Jymi1JmsWcTaZi3YKHdGaLL
fkzWRe0QhRIACqGSfevuqlyGtMfglBbwhaCXbYBUQsVGE0AUSfj6mqjJGBdVltbR
13HF0Rdq2alwfFXeorS0LmQQZBIY/HyHs8oAN+Zac48IDM6VJlbn7NqRex4/tg9U
tvBLpgGBEbKcsawAb3letbZditxuD/nc8ffFjqWRSZ23F5DMWXh/mun+n+/WPtcD
HL+SqXp13SkC/tOP8SatI8RZi71ywDy9WUJ6EZHZ8sPUkB9BfI+0usHtuayLtXqU
0ql+knctn335NZ02vt9vCYxxwSxMS9eYQITxT4kyRj18mSdiGV2yhHHUHDZmYVql
B6bzbSMKhFsDvj1YJ0lswJKYaiECy+KcFA7IqMPuxKUCP0VMbhtUP0IvUMv75OTM
eOFO2y4r46vI/yhInj7PBsp692ZIW/Z5iLh6Wa+Wqgjzgru3xqUoSLUAt38xv20+
NvyAX47msvLedwSGNn71RafCaqrViKhZ+O6QvA3zQCDMWd36ixcL1bcSI7Q7oW9N
SUGhe1AAdDOJxDNbZPB/6p0K3mfgE6W2v84AinrVNLNyYreq8touiOWjgJFcCX0O
wW+Ag71BkP4f1ep53QH+VsXJ4krK2YmENQfK5OBFvQFhkqmGpyupi47UST0mEV7R
1PzWE4/WUUR1CF3pH/HmcPIXSfpD2b44o6HmsZqIGTe+wjRC/VBMakDaUf3kgedK
2XTIYmn8UH4foLLqR+qWxwNseaTQBEyAHOU8lHhSJuKADXs8nXQrZMwIHX95h9Bn
LW+Vrqpe/5QI+91XAyrZfq90CCfr6tGRm0O6pIRa5MTKrlKo4zQH5CyPmmO1GgAM
/HokxDqg91dR3sY3SW5HGZIAFALIGkNf4pgCr6uixWAWI+58wrz744Qs88eFIMp0
r+6f0IKb2vnhUxJTaUJJhZXpcVvWd9TWFW6O2VIyzd5ltDw3FPK+zVoiYge2SPxa
MDrPTiRF9HNzMWwImgw9lRdMvXMKeFsgThogrLs0RR7OUOtISB9etOi0J/VijPy4
IGys4R1z1apuNmIGXeRo84/4WeKJYnNPRXjSMt1YQZMyXa0GhwimfmstrGMIMaf+
PIo8lpdNTmyEXUOqVaAMNKE4TU652NQJBdCaxSFrdcxeJI1FDX4OgBSGGOhBstoV
3bPZbsiec1+h6NQ0fhGJujG/pNzYk6rTq7ajvmzrlU+9zl2ruBgtxzzB26ooA4uy
1Kq0lnoOjkXZhkgpc1Of45md2rFqNXuodfn2LEGTk3Etm9gkuTfNtk0mxbi6xBMg
nm9kLsZSKqubuXQVsYj8LfVLxkxHtmU0tXHphspSgk3oJmMhnf1rd0yTS1WBwYJV
GMtBAytEMOQjebQIUaoecZSSlvaFL0ck5J1A7PWN29UagvwHa3KXpFrGODvIuuXN
A1dV75V3yeufCUyNQTvsxptO5NKHW+SaSUtnLuP/Xp8MKrYKqRTf0/+g3SlPZhV9
4b5C+g5NCDybHAkSl2QftbwrxqGvCjssY4e3MVZg8I1BQ6uaRyOohai9ySb0SsH2
sjsHmpqRTRrwAIvg/VDc6LslEyNBA5rZ1ctv56+Cxqagl5P9AsR9Smu66EJ9nOei
uQSii33z3L+r8NfXqPOADfq8reeujZAjIer6Dsib3Rd7oaeKhIqOMcLHGFvS142a
OTGhlQ7EnwE7Na5CCr3nJrT/+/rpkIrVT4eU4hWQYsirk/gv6R8Nv7rZBDjdsHrv
xPG9bMF0fQp/lsAQ3sOeFB+hO4DFFiZa9PyqIUW9FVHf+hHcE7HdJ+TRBihsnIND
NJ8/+RckBco3y+1HpqqZ+SYSXAykKXGEagSQY7rijXbCVkU+Qim7eKWMs8Cy2qOQ
rXQmK5EKx+WLlprYIAer1pbEQK8IWztvVLN9obXOx4+1q1c+mRvEhT7hGDCUHONY
l3m1eitkYITs8LNSdy+xeMjamKsASNv/rX0Gf1gAV9zoOn/HLlYxfPNLkw9HZiPS
HftT7Cg0N8POILfayydpXphZZlPHqNKqjs5CX8nwa4CzlZzzSWIsVo5LczyA0lHe
2MDHolHvoDh8oFDh2IAisAWmA2FR6YGHRLs97y/4uJvA9H879uX6tzI9zGRAonEk
maZsiWZFmABGu8ZA9FDJt2QM6kYwgEKzS8VbvgogESo66XXEq7HP9kH8WPUU54Kk
cuHKnhhSMq8Xh+Vpymx4ytBhl8RCxeisHIP62pHBhtVdok693eODMW1jg53nmXjb
iORXO6XlCzvMHalQBMMClPNIYCWaDzGV7ez/Fe7x6UTOv8yASONgJBw6AyynXLoB
ZkvW8pQRLGKE56TNmUs8qtMIOWGi+h2OsdepTp4aD6RJ4N1P6Kx8Otqh6ExOv68S
DConrZd4SvToWReMN4EW+fhI6qZODm+KIevUtgBrI18QGBA9OjshtrBU8FCP3MCT
u0zkMTnhkrTwzxUVjC7k5RN3usmeQlnJhOQvh1UBp+LjPMxlx0YCrTRn0UAXXyvE
lenQlH8yyiAHCZLpjmwhZnGVSA205n2ME4uzZdOTOH/4/iCXZNYm+WQetLLeHfDN
JcwHKPwV+fceIN6PQUAcrguG/dSxJ8PZzgEX6kv+OlxlxnGPPxgRgdeD2DU6h7A/
JVx9+ae+vmAtgjESuCOh8d7wsFKzQIOCAk1tkezmglgwbswpkFPoRr0cse7R9UGK
h1rTRfUA+go41rOxLGIc6YnegTqMkRgAWbu1RdEUmbWP8/Q9K0dH+CklhE6cgRL4
DU0grfy1pZpIOnBi22J+KWCI62o+gyzQKG0gD0gxB4+1hFY1LeW5yIo/De8C6Cnm
VXOv6HLRIvYIkZMDBFb1EMfTGL18IhfADKNyA2omQ4tXg7kgcH36ZQgoFUvKqW/4
bCtyxzVOS9lqd+Ih7F5AzJmuA1GB6swqyhjQ1YZnCbGcKcJCvmmiOXMCe/VTWUuV
ipPUzmpo0bBks88L2ik3XUDvmP8V5qcGYCLEa9i02nhYs+t9H3iHPL5SdMp6w2oh
22RIdH8Nnc2eoFQ/0yiIaMRAoO8Xi+aRCI+0AvGm/pcnWG2B7B86FibestjfwD/l
DISfc0fwFNaHyAE9CQw1xi8vvsaE6QI4gOWL6K+SDH30GfEmPmtGR5pVArbkr/ct
ddOkAvmoSh6i4JMNEi6kiZmFovyB1Ior2AJI7KFnb2PBIGczis3HODtO/PwuOZGW
zgaRmg57peq01KX5UYxdNCv0MVfGdIgSrs0XwS5+jbj+khwHj7ZuETPgr7fSyDAw
07gpINA1W+MeWyvdkWB7Scc4EUiXkaIJW81MVO+7YvFFqOzKeOdJSq4/Jmrzys9M
KgXnbbL9uWTzSz+A4pDYdvk3YCxD4JqFMqj7/NraxUeBBjaWb2HMvVXZT3Mx1S29
1YI5TlQOAfhsONCzjE97YKlLBPNnsytId3jDgbtYeUUtREvbCebtGCWg5EnMqLfg
7fNSegh1ClNQJISSmrI/RkrZlP1ZlIEUc78NiWuro4xYXD3aQD6UsmskaHOuOWrx
t6XlktBA23oVaVBLCqqno7EhGL63kTvYBRWA23YiTTpqb6xHGZY/DJpXj/NfaRBR
DmAzeZiXyWZvFIb99ySW0N6C+j9K486p9ZU78Im7BCz8WiWKkHlpRDKquLtgMFVJ
hEXQMsggTmlE98VpnGPF1DzOaApE83oC2AN5qkmcrFU0rd7xPtJUrw8CCtt2PJVd
8++MDDCJ2MacXE5n8sGHpps38cItueRyBOtKQWDgQ2hYZL2e44zxkzx5hsAsDS05
H6yyMazUByouVCyKlmAMXdtaWSka/DLstoBI3MZmaIj4vTLhpnfxbxP+2JoDHp4g
3xuMv0cpisOeUHBk3iQclD6SNoxb0+lVTV8cJwLtYCpNsJwdek/LGpK0+nHNa7u1
libipVMqwmguh2IfrxHrOkhKd4VZhz+S7nx+qYPBxQkXp0Hhq6DC0TbsktVyKvu7
9IURFwHpOlVauZ5DVVilyNJpHDJn4KVxzwQDfVFZpsSIgPj9SUZyUfFw1xrS9Hdg
lc3S/N6d54oMDB+kMvNWW9P3fC9VVgVewv21AspP+ugohW0oScTTa1lRUCtQHsg0
YL7drN5k0Hyl4bgIWiy/N41K58/2YHKyTt3qX9AKMSbS6Y7dFlNQFX5hXPSCJd3n
Ol4rC7bS446Q2BT/ZiPkYYntkd/LqrKgwP9+sNBg3mEKkpC1vs/TFxNU2orTPuiF
JcUMA6uMzMilSV07ZPONvn8cuMmd+81kjnmP8MTc3jUDuVhG3F02tcw/c8SOiOGU
BBInkVaXCf1GNL7vXG9ge9XfMy7nP+KsGwGWvCX0ru9Ee9FVJ15idp+L/7iOBRPz
PoGgvf3WVXrhGvkcOZp577+pq6kzDO+OBkMq0flUb48I4B3Qv92fIX4EAEctgMCa
KXreHH5AvNBEfe5oK9qAHbadfEb8O8ZEBuP5e100NEHWc1vTsTHZ585rnkG0V3pP
OYFjNk/emzuHuYGvEeS0RDPGHi87IkPJBYRSXr6JoDeBid3+u1xvQuQbjetZ6EnS
LbgTLVX3r9KTjHGU4RXzemVKP4/j8chkI7GEl4wcce6ElkxBhiBXjqFakBJE8yF9
H/LyaV+IiKiHdVndiF/tWIO+fTu+SPH275allSZqz2VEbjvPx6Wy6+6pB2w6l29k
9oJSumncl0HwIrQfQpM96WBzwClzVRnYyoC4SZT9xomabVtlaCTjbqDRE3Tlksa+
QrtmqR/iSAt62Bwou7Z52EqKAV2/3EJ9pUidewir38H+LJgG5EQ+x2ISY04+jrmq
Ow6sVs0Bi49ASYNFr1B3Tz4cHqAPTw5p++1c3pyF7Q0v8rQNFlHB/xgH+s8JOF7H
1scrqd3FsGGMha1YyOKqjeoIi+op0Xehh/vv7Ea23OM4pe5znK0yku6Vl9626DHz
e6r6OHdyiEWrunfgjX0/OouZni+EacpmdAioc/mKgIfSr74KOFqx1shsXo2g4WYu
De19nlMHzwMEbPlBWzI0PZJ0AqxtjZRM404FUR5XzixxPfFWJfFKf88SXeT9iDop
7lIrg4pq2jdZxy5RzpVxfpUlC1NPqlwLUAu8E07AO3wKwImOmTAWgWhevxEm+FeD
NDxpA9alZK7yol1xDmf5elsPjvbLSjWUJOO58kurprF1w38s2ljCFD/TEMMNUbbo
Ee1EyOHtf80rVaUb/W1PcRiizRPr62SyUT8yE+A5gc30Fui/uiAnREm/Y0B1m4tp
haFQ8ZWiSwqPv9bARNRXY1LS17/UI4VzIJ0gtoejN6dhuUUtdNaDs/TfqaqaRU3E
gL6/6blS8YtReT7koKTriwqlIiczuL7kshvxq6NmHmqu5bJA6S6z8yZN7Zi4pZrf
71krL7vfZ326FxC2ZcRULMrXB/E6NrOenCOTdmLUQNpRdfJ/OFCQPQp4htr8Oq/U
/ARDipAubKpHZLrBfZKUmxfygNKvIQ4CBaXmRIMvYdUZXIx5jCh2+yqxhujxz6d5
mUynw/qWMMmc/OoxaUYXSZlbT4TXuvM9GmdGnDzo0FPHEkq4goxmRkjylf1IMuED
Tk/OcexAgXX3+ulUpTwHsFv95AE4MQPDEHEnbDcySFrhydb1QGIl0eg+TIJcseg4
mM+Q3npT+jzFQ04no6Cg/W/bby1RecT+9TjbZm0nY8eSX+YAXH0S85iUbVJexWNx
4l+gaH4ez0Xy5SZeuE28zu71PWLEJYGECEuIaxwfyUdJMHkWSrIWEFniWEqGKI5Y
Ov7Mmx4IkeX7LDWVfWfeHbi+g+sxcBAgayPEP/YSMzDg1IkefADaCFfcLMdbtzwb
19LBRIlDSytgKK3AUepvZV1UPQuALYzJ527/r1rQlrdxGZIZ+2PMYKW+r1FmyqOe
SzY2Iq6AK2f+qn7IoT85dd6V31secTX+/gVeIiKSkvqIKVmJV3IgMerTPAOIclGf
XeM1VSAzO+DGnNLrz3RdXCE4rRWq4sxHxecgDGSJ/KlsxoiLGl4gWzIGMNBXkJI9
3NOwPOoyzY4hJVbS7Fl8QS7/twaxm0pksUwRYZd3gM2nVM741PQtKcAvKx0ZxWRg
Uo2tdwmO0AHuqj8u7gteOyzEZxCrWVCVyeHfXzuBfI5o6/DDU5FKxh16LIJ1tQ+K
eehvAxMq1I4AwgcFfn9TBjFDWHNWeaZaU9ooEw9yzgO9BHanfwkuQwmsUAbR1/qM
KgWVsBBN3Cd90acwXwb53RwCl4kZe0TlloUCPLdU9s4gvfVOqftva07WedPdAGLQ
o3w84rnIYWJLlLd3Aog6WwoTcEf+DjfI8x8pCsZ5dWtrG/wd+N3i4XIfyMVXEb3H
n+WRT2ZepjdHVIniy9T7BwzWp78tm1CrVmQIzUNzRXESbHu3Tp7IqYenuLkJq1iT
SLOOg2VKA6a/pUrVyDMKIPHvTFUVgvyidBysLzROpAkxcKmyqujkc3+IZz18IKOp
bx0JJxt+ybiWZZ+8oxUGUZlvBtdQnuyaCGIp02DwaiAaxdfLtulQqodRacMtTYEa
rqIse1H0gnQIfX7kZ9e2FZZblzKWKFb2Ju5oW08S/Wi9cn2rCXA9WM0I8yJwx5Gd
5PoY3NVzjjRmvYEL1GMrRxtHG8ijIkMs5UgMP7RUSkTl41ejj5PDEpWTWZl8p6wV
TZIhGavhg2tOUC5XmEx3gzxSKoLgl0S5FN8x345EG90fPzj3lVXb7xggPFlxs5HO
ZKp8BEQmuXlqOogP5hEIbP5Ed/ELHxSkrox77uiXOZAthFkr6gCgiRMPl+n68YUZ
DYnJRbe/es5oz1FTklQUTRv13inbJzvWEAgO4fODFqqnRpAUuZGBk+SC+CC7ynKc
pMFaew+eJi+P517KdIEItekucMqF+XlzIPlAAma0ZhjwvojLdbOCodQFq2peRh7v
IUxK+jbvFLDU1ktRVD6xx2+/3PTRm93csTDnlrN/2RyHMAaWXXjnWllKMj5c0u4X
zmmmaYA4pYZIrRToPRrbY0j/pwxCw3QwP0R4/hauJr5fNPhyTiot76Xp0R8H4fIf
/DiUmMZYrpLKxrFBTI0BpbCf3EnV9L5UycECnJksw39EJ6OKnnddeHcHo93vexoI
sAYcZDHoJ78r4wtmw/RO/CAJ6ups6BdaNXiwxjoag3ETb7eRzhcsPM7uYCrvRAdV
Rg3czL30NjdpfbOX9HGCbCLuGmhGxeohuC4k63M+NExyVUeTRVAaLjULcjCiZDKE
lNkjJ+/8380aG7uX3jtTb3XrQ1G6ZcxqmW8xI9EbtIscYWmXdMy43elwxeLv9n1+
2iO76TPloHKxRRp3VhCofA3M9GRios0gIc0O+EN0z5Qy07VVhta2zxRuj09qs2Tp
5Z8y50EzZcwHVjSur0KOQkqkxSumiy21/cPhsaI/HdXOLZerOCMkJ91BRRzh9S1S
zBXyXYAcMRKRWuklq4a7csDzj5xOqw3qiiirEfNYRtML/7o9e2M5cEgmkhyjQQ3Y
NUSQzJcNkenwASl2ziH9bVYq+izh+iHj47K0kRYfLt2Csgn33/1icbP2A0XUR9iS
71jKRPEnJ7gE5dvoBvpT6YBrhGXZOEGywrFaIB7enQr8OIWdbvIhoQanINpzhTRX
dGKnrz9lDDRlXtaGbR07yZ8Oorf7uQXGTxngRBHSEvoeRNJGc3G+iwE73cwZIfVr
mR9H+Y5cQyblhw/yhH9FUMPE1lDTHIX8Bwyddc9P0hom9ePgsT7WO6egu0zdhl7y
WCIyoH2SJgFVXjrd9PAA2usp2ypjJTY++tpzOu90e0CE1mSaTNha6/9nfhsGj0gP
Ev1Xq6J4oG0Js2qLqryRZuU2GIVRIKF/VwN1rN7uRvx26MH55qFarbWQ0xyH/NRr
KU/NfOyrkLLDujXhTemLvlv4LizVojhlkeaAjBEJXZj3V4C2B5RvD608HTht950s
wk38w93bHVc9rHR3cz321VOeXK8pSR5kUljZqooPJSE8/4fXsLDEzBUR4ArzPohe
lAfjp5HE33Gi6vAOv8byydasJPPOA0YtS5sfsAgcNSsAHfcDanx7kNKK4PrFzBaI
9F+6IIfwFcbU2x7TYmGTPnfnQ6RTEw+9Kx4LX1LVTO9cO0Lr5VyQLG6atMiC8ibs
i+mskKJx5BjiRreDXsjnYEQQvT18gd5rusTd0WC+517xHplfQVQrOnPzgmjwRTzd
XbOOTbZzKrX1jkpKKVz3XD+LkUWuD6h3UOv9qY+Rm8wS29QScpFf9f6ITkKJ8pcX
IQCOABjeIUsuQOKqFPptTnzybce0xoFOUssPpMCemwfHLA3HQACG+xAMt9nJ2SUE
A6n6KSv7LcBUmUQxUBw41adUM27XBN1/P3AEnPxMti8ZkMRLtac2jyYbyPUgnqpW
XXyJ/KEL0S/kJZrN3Aah1uHeUM6hiH630E+MHjDOksk2RwMdkI8eZWwRyvMqCh/B
OvTZOqui2bnvAbAgb3nW7XfSxf9G3ya+Wy3WQHtGfg5LiURhHcKYqulosu07gRhC
sJyXTeyBUo6i5IorlsH2ddLR+BJ9/KvFN9LY+9CeGTZjE2eyYPSPN691yxSJkIq+
nIIjFScTQjpANo3Rbiq4wglw+sRyEed3fkDNpaemodd6SjlsZt3PNrj1BtOgqrXZ
0g1EVEaYP/wTyEXV9/gz1sHuXlaZi0p0590mfSaUQuMm/iLXYPmIKRKRXHRnDXMq
/OxeGmrODaZ9eIGB0HsfrdVMurwDgAUy5vhBlL8CN8j8Kl6RONNbR95g/DgOWlPM
1v0jcr/yvKQe8HJc/QcSfnojx8S0hAfYlpNouEySxMU6ykWA4E9jshrd/+MjX0qM
QL+cTyAVoTCSGolvRrK+nVDElBJHc+oYk2pQ5r0HutEcTdA7nBiqy5wggFZstYfl
kfzisG/A0+xqhlm+aL8uvjGN+C6mDfrP5Egur2fB5mtu5x1k4nHnVdXoSHNwCRQU
evBG847CfkrtIQgKjlE5A4MIR6gI2YoDQAIMXqTGErEnRZ+VaGnR9b18T2fGv5ep
qf8HVgfrucIHKK3h5V9I384UEsq5+2MOFGIleWVj/vgFDBdoQJk07GcoMy/O1uWJ
iKugqELYy1HpTJ54Y2BOGSrUE+eP1NFkkq8uBQr13rAi5wiuXg+AOAuOdMcWKCYw
GvA0nZff7OC6F6bfKLYFfIPFjgl+o80p5mJ7oBdulay4xhR79JPV9BOvtvLv0J4L
2TwtvpXplefBGB77nPI20xAu7uu5aPT1cIlQMJ7FUENf1YYYXgNffWP3aXjj+HsT
PYSDdgfiymTKblm8U4wqnXB3Q7Su40KZVBKjpG4aID0on0OmPbqaRXZ1aJCrxWyA
erGv2+yZHfCdM/rZ9R4FOeAoeBEx0E34Jh1Q1uiNLrLeIUyBKNpp9Va4eStWHTqI
KGssmy535jHlKIr8x+iwRo2jA+0BuzEb7nQz4QonVCE6gx+P8JWXucWICtzFUDJ9
Y6BfoU7w6FFQoJS49DGMBv8f+onPzmRQiVgLVbJhY/7zivc4pbNSQ17DJ7JStfLZ
0bZUduv2Vtx+pCIAUn4e9zd3gH/aUJnmPNm1kjXK73XhjEfDXTaCeJrGls37iuZo
fiL6SOZKkGJRnSLbr5ihX9rIcOuiwncPcakxEkxAAeBFcPOG1F2+Lb+eiQHFjLqs
dONhfV2q+/LIpXrG0UF0wzYFWbtyBLX4XYh6J0kGUqY99zYWOE8FvJD7En49UDVW
9RK97F6XbPso5UsJYywTueN40ctLtaCIGd7asPFqeS9/D0TzJdxjsM3A+i4U0ixx
aDBeA7VS/XGo65/BR0oRzuMAC3eW9bIhWRJAfPEUnN2bPs8VlgqEIcJgqmH6933d
d5zKMeypMMXAtVPqrKQZVc/TVJhfrOc2tdQLowhtw5QfqraXppJXQwe+682t3xkG
TZV1IKwl7xtAyi9uisEZBqLayGFJ6Ovwfz+SgyPo+sHeC8ugl0GDIXwWSHsawQC5
kZUaQVhq8ObKx5URu6F3kixz2IddhPwHLxEesulh6OhnDHB1Xyii5UdNsl0bI7VK
QL1jbMCg3eOQEZiifU29xQhzmt5J987VJjUViTng0jG+j/QiOK9Z3ofh2cJ9+acI
/evoJSKYpdv/lZHKmREVfV0cI8QD5QLoJf3FrFeddN2UyJ4Ozvz40J9rFiRZQSIw
ejLPX05hOtQ5RuVXMzUOrWsK1od+ar/OsOenvTPF3TL3RI/rSTYwjSNcIqhCbK2W
Yb6qygpLUXe2zkegY9/rfG4Rc16o7cKnkEBTZLk3z5f30PYIZRq6Vxw8867T2as/
PyGhVCFAADnAUrm03VI0WhU5goPA4Xi+It7+XraJrhUNUeO/66h3ebeMmq9ylAHo
QHyfELbaW7bpe+vftIWmtNAHpYTMysOmoZa6G+m4jc77vr6FIl44AgwqRGR/qY39
QOF8T2sjM79AYQ3SAqQAT5OHUhwGafVzIoJcU+qJByH6RgsMbxI9hWq9hSvz18/2
sQOHO4w7HrkG452/YQWjZHHS8dSGZ+74vjhyq9lxB1+XyI0YwbTWQfFWMxeAbABx
wpniIGSn78IH/fBo0RyJokusc8XuQTM6QvlYcJ3+4kqCpqXxuXdKU+OsxfZH2JQj
tjorACXWwzNd9QZQNmO/KEX5EQrkveaOUCrmX2kEi22/0+hyx7LQU+z3MbQL2YpD
UYlqGCLbBrTTnhMpR9gEeXlYMeMfvu52DQ7O5PIfmyBBOYshbIl7EnF45Ju2333O
tWF4gbxhJgZC9x4GjvVeQnCrg39P/ylmHK5Z23/VfXqEk9OoxnqotS17j5W/Hqsw
EDAv2yJzmv3bzGE86x3xMS3ktrYSX1H0FR/k5jKhOvSiEFpNv/2hxAH4KsibSuoA
tua1hRX+uuUHM0OGIh3fbQ9xGLFMDWoVsOjOmXoJGCc0OrJkCev2zlNSOEZJTlXM
S/s5SnR/qLOqfPaU83TEauWPOxaAmalHjFfDLdzCUAtWp3hnUC0BpjVIV2UzVeLm
MkeJHafQUMu5JSmpJasgO8Yvhp0iAk9QhJjMopQVwoARsUd5F950/guqhXOB+KOc
QCeFXa4HU7ioz98CiB4XJCoBBoTf60PvIt/079IbahjCzGi4+mawYN+CDG0CTelY
yDgh4vMqt+AiHRfXB2Qne03I9W1PUa/hbhpGkETs9SJ6PsYZ11LPmTLM3eFD11VK
EdSQYfemn9lHNVO5N5wMh5BqTwnFhNbUYX9++BVVVElz7wEolTZZ8ZuBU11a8MXP
jvVJiIXhVDgDd91YEmT3ORyP8qQ9erIXJajo9had+IJSA6rXtQIx8XYGxfb361jI
FxDbWUt5RwfDM98fiJmlK8WnysbbFuH9fif4UKAWKzdO47D8mHr1oeIeTZMGaLno
f0hIHUAK64mloLtywA2whyqDpJNI5pZU6jtuXwMR/8x4hlYfpAMyWFpEzIAAL6OS
RL9RbrSUNpI6uV4pwVeqYCcGXdZau9lyWkAQ+dWDNlzEKHzT9Es3iUGpmv54vKGL
GFNfY90ABKMZ3kfET3rak5PGFYaEzf7Bgf0j/WEFvhTwYutfH/xrNG4OAYi7Pft0
mlBcZghSqmKbkJMk9ja/1w8ShM32LAkupqiOGM0IM85U0wL3cY8WZl4FB+O1luLz
eMYApCWLyRZwvHsBv1qgO6+BhVM0L66anuUPgK1fcXA8RlKOWwyD3jHcg3lyS3cd
blEi/P0q+Q5ii55qUJAW3qKBBGvDcxy2JqZO2AB1l9pb9R2DwAdioG/YLsPLUgY8
pGa9Cs2vlGDX30mucbqYmft78iHwztQGaGA1mLRXv2lJp7gTB/GVeC5pAaIuOE8g
5y83M+ucbu0un19nL9DbKAK/vUwdNBB//OO88o9x97VIYnnah3QSInfMyBU7wNqz
w/F8tspd5irbPbtTzKavXmxBvlIYknqu+HcHoX9dG6eXXqbawCiMBySPgMkqrS1c
wLgd8qiPXChkckBy3Qgw2VfQiM6l8+xJ3LsKJNr2eXhdv/HvwmFMm63lSvVZwJlA
BfRqXv2PnLNsBsVKsdKMP8aTn7yKAhyVFI+1FZkq67dCgnf4MGmwf2TqEMKF5tII
po4Zo41tJWhbsbN1zOV9RcBYRbu8Czp9/nprCyooN2sSVF8CfFlQPdD3AxFaAp+W
gdk7gfBUO28SzqQm/R4EHpDLHOlcNwXxcLVF3eO3oJfmCa3luT31eUyUHB3OkZmN
+7WQUTBrHuKannTsbnP5S6bLAoe6FPvZvXgFm3CtBmhn091adSD5+o3uE6TZ4pBP
rCp/hEVbfE/WxaZtgbpazPPdUZew0ndBBEzyJUHy58R3wJ+Eh4l2PUanVxDT+UDQ
4htrlwINSgmQO20xz30UjGKJeadIt69EAT4i+Flibae93WQPnKiBPUxI/KDXdHW6
SoQ5QlRIzItXZh/67X2LV93Xrdt0shPdnr0OI8+7iGiDoHvXL7hxgqWifXMvQwNP
KW3lqnNbOL9Tzdd6DpaEmn4cr7jAiWDBfJSPa+TNNOVsRAZwNBmuHnICAM/oz+EB
D+9oNaMWpj5+y6xEgwrbXweRFeVXi3Hj8FL/Mp5hjQ7JM5HYDx0ZHs5m2nPf5eyD
LjcLUZzKZb2wuurGopvUtQIjVaIMCQxsxvGvz+rjjHo3Y3NgHfFrYGPHn+lIsGVV
zL+dCYQOsCbu9JWlvnqooHiJ6q3VZKpOhQHRCH0ywiZeZysSXJE4Vsz6I+s5Phlk
/TsLgaW44LiHEbrsGvlO0gZG24/J0dBjxgdAOVO4wOtwhHHTBcG+hO4I4MEmJWic
DnfVutjUq4CE/pNCieMQPQc+5ozHsditw9KyUubX2H1lGTJZd6h1UXRwF509lWBB
CZu86w56iyNVbQoh1+ssx0tukV+9+5cVGh+VLT2Vkg2nHNHBGyIwVJpmsGh4y4mM
2I4XEcoPfvbwhBcxda6RG6CfOXUXV2BG2a6KCRhRr4e425W7YyJflNEuv09TESMm
7GJwbUGsJbxRKPCmeCJk1hlhqjaLYkD5HWYyLSXK1Cuw4wpHiaUmyXa/0ha8sLPz
z/zUiVmyoJx7wgXm9rhBBmCBtegzvFOPCdLkeh1RdDLEYBucWBo1kOfDXfo/KpxW
drGkK0/lrA6/FsknERlmedvZ3Iwa0pUvc2rgTNgU4fwGBRoExsO+jdeTEA6EpINV
nHW8xk3d8Ymfv+GaQrqOP761iVOeeX9Ztjj85g0Sd1geAiU7JWD9yJusTw3iNlhV
ivec5JZ6xjPQQrQduY7L2LqBUdQT6qXIcavp+HyVpmdJS/ArG9WBazUMbkBOoK3o
uifU5Hsn6g+WL0Swwf9Yg4gZg+GaCLeKtUlSwEQzKvlOcc4UkxyATuRjVZiuwwoL
Tg23CBtThcoNztvK4LGE8MucQQAFiSpUB/sMb5oyf9icKAaXqjoPEfI37T3bNi49
g7cIYkz8vFj93VgsZgESNcMiV6Lc/HaqOcejktaKB7pV8BKyiv2HV7QW4xc7vwnc
9l/MlroACZjy0X/bi2kFBvUiZ0zmuQKGLYxTwQCIAnK6NsR9ro3vj3z7NNwHZwDY
uZYopqHG8cHYDpsnGWMy7suhrqjFfESLhmMVzAP4ao4193BkAfInnpIragw3LpXT
YKxOaMjHQih6q/OrLK6ew58TapUqwbllDI3mfoStdGqDDDNkxk7UMHqsTzbQhrOT
9KFvDqJm9kpz+O+Wy9FxQ9OhwuIAk2dLAw8SLF7iQ9f+EVKdtRuFICvt8aVgRcoJ
2iugwazo2NldsniqYSBQYY+vrknSIunxsurgmqdVRvbREPHCzp3Lp0PogWd2SHxu
iwsHncD6iF5MWyT2sd9Lkrqypz4KrWIl2tulVNcAnntNKTHw0+biXwmL0Gtw9DnT
cRvsXXKAVIM4Eo6GQjmJoYtqD1stYNkDPNn26zRbpxpguK570KbZjs4bTfOM5hki
RwMBgn4SgOHhWxn4pZAGWU3mdBP4Vmwsbs5PHxQxjVgChNCLDxhhC8fiBBr3D8zd
nrgdy8sbBR3RQkLHZ09T2X+EmvC9GW1rh/EJwt0zsk8+BLlKno9Ql76TfbWmskow
KqQaLZAoi5j0u54mJBmHzJ93N6H/OjZIxGK9gLaxBaxStnjvoWXVC/4KjQdO3nXs
Te30TtBGhgdz83cHtKl3QAFqDsgsfNrWR5xoeIk0kKa+C/eNuauYm0v7lRupbdwi
xdaovZi2lwvtaA7u/OibwDXOHEE5jgFB/CevYj5tPuYu51SqMNJbfHCFZJzS24YW
koNvkCjKoweeq3L7drTQIgiRN1BTj6f9n8HyacCBLA2FC0TNW2IBQdQgMiLR4cBh
L+kAP5o6wd9lBsx4r8UxM0BUH9l6GSqbEmyDlJKzdPvd/EHUQcXru8StEmb2Hq/+
gqkwMk8lET87pCv7jGzQ/HaFmUVPDf729Erm3xJZoY5xuiHRJdvn78K6PWtugvTt
IVu6OyQCCFB2oYkZBzIMdN9OSqNepi7HEWOCDC7KO2i7NfAcCoa9QuUUJlUpp0ho
DdizOt0ZwnXLV1BJXg6TqRRSqb5Ix9V5pFS0FWOLZLXFAk9yeiI/ZMOHurHtcXkK
uMQDtsDmOCA6FJcF2tfx/IvQAgCUHuwUAOPc+SCj6POhFD26ZbEw7zk9dT+FiM+U
SFyDnpCaYqeUuukpqBtAxwmckbxAO2SsHbYpSpMMdhmVIAU2NgFFioLjQC/3iH+z
hRkUuYELICvNSbfnKU/r2sONmHp0s23qZwG1krbN8A0g0kztMEvza89kE0Q5Gr8M
/9vB3maZzKat8JRi83ciQjwhJTi7/RrDkdzgSCp9VeKXn0xdzIzsC60gsetQLq+5
W6tdDxrrVqBCCH43AV3zJUiQzbtB6QeHhl/2h4UstBRZrvcIJ3awE59Ptsc1kzg0
pi/39FPqpcuyK6LzKcsOcISi3+0pCmde0ZijhICpcVZ0iP1t4RKGH2fL3J9BbehW
hgAJlD6jgPoV+2deIDTgTeXUi6x3bbYrWPtoKar96f43xPDDaPehyE0m4SA3xbrR
Xo694oqfaKAzUDcuqHOTVWgIoNS+BwN2AIa3G2cxwcXDFfRprLnRHPByxlKg0bHe
wyLdRn1y9FoaaRFVjcShwJnJJBCVySyDdSPWTsDP/0V8nqQrIIptw5QBAIrOotiD
PtUzXMBsq7+EglPejvXNeqr6iYaNJ6dCn+VexXNKlV5KVySCx27VT/Mz6Ykn3s1t
3sF1awu9p5uyEgzuuTfP0SnZecb3JlwQQ7goDb/BzS9+AEQPwowjz1qGcPi0aL0W
ZdtGzKsg3AsrdhWFQ7krrzF+QDWLAROLQK13pGH7rUuyRK01mcb5OT58j7lE8e+l
HfiKBoF0x4g4HQe0gV8eyC86aWSsNaHkhKhdUi6djgPLGPD39P2Y5EN7tp+HUdoq
8sNovg0QYvA1FkKBE6VLqKtgZIlhDOHFhzf2DYCeYx0fOMTRho3yhjaKq7P9jWhX
YACsRXdhTksxbAPG67J/euFPsNfvLmy+hBKNfR8AWhPAeyq228ogo7/sTG2t6EuJ
gYkjkzvHTxqu6UUuQijJmPNd3UDSpcRIupgjOlOU4kCFEciQYe0pWj7RmbGnzL9+
YM5GXyOhxKzkibC1jmjJFQcddQCJZo2NXO9FqgxKtD0KIcpW187yIM4Ag5Ip4bBq
hHJeTymqhBwKmqI0OO2fJ+kpTqJ5I1zFVoEJkQj3rqwkvdhph/fiqI78wDZDse/h
hV3BbARuTokMkO8T5VreP79oiJrrCnmnTK0AtpLi+K9jKTLLJxOOJj5kqGdik7FB
SfzvYN1mGe8TnZXahwVBz2qwtK6hqL1g9aOEMC7NWVilP4pxrk2ghzAYGPBKJ2hu
v7CCxBRIQQAO1GMxUhhmybOcPggzZdT8u7cNYsUoFZsDJQ2Lqn42+a7zE9br+FCR
iKkvTC3DsD7xI2AsZBMemLR7UXjLrS9M1YwQMwjWLeQG91CNWbUNX6EMyZA4+lU6
2r+jYfNfcyVHzECTDSpfni31JgPH5uSTgRsqAc4dCqm/PRSK01iir8m/xWKoWrQ8
GOERZvzYFkZJI2dIWnS/YpAe4b9OWZmbe0cPv3l665J0jnn2allimmfz/0+ov+Wg
cKviFx9fDt/j6g7dlmGDnPjZIfBVeqE0sif0t9X63k9AMFcWQ6E3UDlMpCvH7FzW
lUrS4ma7ZtJ3UgmPam87LBhV7WBFuDm2FnO3Lq85S8keLeJY+BAgM/DT5YHDwZcY
BoYxg/felvJPUqnsP2bw5AgLhAWeIm3ROyGCO/LcM+wo+BulxqibIQ+t29PdKbA+
XD+zKudxnwm1b1WkHExm2FTuBUg+3C3MLFNIyu+awRpvSU6IP6ZoazuQhI1QUXkk
YzGJLRj8quLdnwULQEu1P7sP4rno7NjFsIfhrs9Bn//VaZJK3z7sXKeU9Y8J51g2
pFgp3+BkhGDszcjWFCMPYayhw6mPw7+KzrzDCSVgZuOle+ntXdx33FB/11ORCaq3
GsGelne27GL5HIgIMq5UkO7AP+DHdqmPg5oVAyISXRn8Y0q6q/iwNtEJONExN+SF
+HccUqgrk4t9Umi7GWYD25k870mkjplxKPAHcDKyGr6Ny88/iNDrKmaQro3AHVH+
E9cUUh6nNbUp8hY0wrw4JwzV6rzpzsPT7rX5MQin1Fzxa+mUL3cc2ra5R3VuxfeE
P9MMH7cjsooyjKZPjrOF8lKVOaIxeU99j8aa9N8J759E5zw5tnwCywuQI+sBYM1I
alT/7DSXbD5/Q1LDkBAfTfD3tVS47nkxPxsW0iFJtB/98m8uCLEoWV4NiDs8+/Yu
YcWtGAo2BwBmWUSZaDEjfEt2buzuDWmMF0LGOp0vw6Zuteztx9XxdPiTGFYlovPC
DFwwATnFr1yAIU4JjgMmvvCYa2ktJR1fnFpNzA/8VTYLjECCYdQQUNyUauSdc4F8
g+Vn7fSCO0dMssaLK9M6xub/t0HUrfUQUcF8dabcHPBrcDM6YbhJOHPfwxIvEoN9
sg92A+bCpLCW4jShqwdHPUy8XoNMRnRyWXai9Ian+P1f2/9uVivFE5SEQp4bWA7H
LNYkhuEukPE67aaGgiQN5ITZYHFogp/QWZtKy4bJ4V2warMqg8dwai8QM/4zfVy/
hUBOkgHLZC9rLhb/fvT8A3tvJcI9xTR23rweREHO6pWHhGTzhRmYBj2mQcP0LgNH
zTk44X8j8I8iCPkoU7knit9phw0t49Rh2NV6l8Dnn6x0qRoleqznzj+/x1V79hJ7
JwQOtJ+X6cDhYdUY7kli6tyHrr4bbw79q3vYeOOL8EuAWtzGc4nY3eV7VtDVQuIr
DdJo54d6+QrFI3HbXPIkwLzCQmsnauAvNj8g0UZVYc0brhBPYwA4QuWv7lNvZU5S
QYYBi24ykrT4FHiSw76tBWJX3W2iDTzz5Awx6cFsEKhcQH7ijIh2z8eeJqqbuy/2
oCcdylERc3azMtHVS4BB+8gM5qRFJBq6WZVnht7cAWWFoxStWD7Rer4MGXmVz0gy
znO3SAVvun+N6+1MWeP7uuIHjoxuH265avDcEa0uE/cjGy47oCBTZ1DQmQAYe18P
TMuYUcGVilhmWq/M8BzxYQm+rHT74X7nWMgAp3vPvOfYK9K/SeuZkrpiMEad22N1
F4iV7bm2bANcin24cccaJfB2DT5oBskGbMsQC7O0Vm/nHpOJim1MtEkUzHUiwJcQ
HdlM/H83fyvA18OlfBNo1vsXhwAwMFy6K2aw/PKacfHZZZd5nWys87WKmLJwIcia
wZjzJA9bXEPSfmruBjdBa6HRm0fk5zzI0VBrNP5T2UsmrZdkkO1ClpkgXJJAotys
lrX7pGfwROIzJkDgUCT9Xn+r8T9E2YF+55cbN5ywqM8ULXPy/WMSXwtt8SMUnvI+
fXD5dxVCrQEmomlFNJDJr/FXLvMgOpZzRGo09pmcPKeinPlMiDO6EMuA+Rt16OhW
dojcrq2YACSsINT63WZZmccmlqTazm+Fw/SoswOIyCDDIDzLN4S0gPAN2PUYsZu1
Uu06ghxi6iJ3MI28MMKyyVQO4qYDhOL4bilnQ6Migvoz/OgcVuzvptX8xIvmfb3z
vCYR0gyvhljZGQ/OX6KyZg8O8exc5jZz/DinfmG8ezR7hAjopc/HFiI07V5IuZK1
WpCuQax3GqTZp+k89yq7SvM/+YJnodi3eNjHe9ezl6SbmFWqp59F9A4uioETE3Oa
5F7LcDmm2aS+HrBKuNOYlhWOro1ffOMeOTT7HHjXyIwr3zm6Ub7KaJrvj0FHOw7i
w+nddRZ18f1PM0QIA9ntbAWis/O3WeZKZAIXuOfkGrGYr5y316eD4l/oVVgLmJog
mVN39/nmlbyccYlMWV/EKYWJaVV57KYTE7/ekTvp3UrPqmpLKAMJRZ1XGrO+io1s
Ie2kgu7kn9N2pYzhY4OO8kWCSFzfBh1FcRSydnr5KdDSwTEcBVL/emo0kmz3rjYy
RSsjAiNXFIUf9obQt5K/YlJGI4esMpWlkYgppIPoL52dgMbpWkW1zwdMMG1/E8db
HgOS352sYa8GAJQKpVB2w7U3hISp/PqlGiQj/v9EsrXmbgLpS98MJCHjgbPXP7Az
sDOfmAZt2tl5H7FOFVyxS5XCIKfDT0p69+ZM6QZkI+ylkykD1rgmHYzGM+7+kzP5
DCkkxOtFiBWwg8MKEwIsBN+z9U6q4Mz9LDanSuOKWkkfYQ9suJ/BGFIBFTTLr3V0
s25whtoRQJw322DRVvgWbT8nYkNUxh5I2CNx69C8xDut7L98NhFwHA9snyYD6cdW
RzIN1ccJa0OVwWLoCR2CAzi6IAl29Fus2RtO3iq5mBYoIHxLgdigUthjsiQ++SGF
`pragma protect end_protected
