// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:42 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c1uXJHcFfOEf/Cts3RLL326RRzkB7Sw9RMoyBeGniHfgSuzOR3dLC9iwmDHEohFq
qDXz1IBoZemkRY1jC9qGBf3ScITOM4OoN3H3a7aSnWQ/k81dkttrIwyKNCT/KWXL
bhlFdjcKeQSezZi26e1RWjUR/G6U6pcovY5hKvpX6qQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22256)
I+PsyppN7VdSc0TGde/fugjdjBK2lhJiWDy0Sg/CELhDGl6y1ir7ilGrH5TnBClZ
piJ5qq+2D1etks5pMb0EU8SNgy1L1fhRr6TbKKa4RwJur1Yzd5Jl78qQOyW85Crs
sFtQPlUsjkhhmBP67mcZmIPNie1cAC6tiKbye/bCAj/Em+d3k55PIfQ1EqlzbW4k
LyzL5IcT6P7cCvTcOB9QSayLve8FhU1sDpJ5dJTJ+6JWQKrhVwiJvagumdlCU7q0
GDsj889fCYibjt36AuP2mHXFW/7viOjVjuZ82sSHn+DWIPj7aC17/s7F0k1XRiMH
gc+hA8tKWhErSi5uzZPBUAlvl+YkpCd2BXiCQYEnX98R0Dsr5q/n1y+FRa7vmvL3
yFoIvFoykGKUKLLAzSOZ1PxcnrCb8f2awhv3kjfPeFkDz7kmzAbOOBuavmvGG65G
t9qhHLZ36Okc6D62a4NMOh71EfmPnAxRmDkPMJhra41iNU0iroD9SNniVu3BuxNY
+dl5i+tojft1PrNxH/RDVwCesyauVVmi2ZnmHh6iREb14qGlmp3lFOIPZIUlq39S
lGeoq4YpdOsPvn5Jue+KothH3ti2Z/M48yVkJffmnL2WcV4KdNIjfg1wra639K3/
rnvIDx6Mi5HzdveE4dyq8JqHcuNtR/LY4GNvlnS1SXQ+COJUG9I0Q/Vebi9gpnL6
/gPEe7WL4SD51gv2/2buvbZ4jUKTKk89nPmwrpd92+bPsAyA4lf7vvJNHtkpx0/5
2qTXrAlR7iIYBaS/evablGDCsJIVRM5pINcLP7A8IUQt2Jfn2MH8A/zZz2LKzDBV
YrKJxk3xv9eNGIZiO8K454vo9RBEvvb2oNxSuIrX50Cf4wcvPDzXz/7n4ILEz4+h
95mkQW1IN4V/2otBslC+PJxtyKP9fB0iGXOpm4wlgGH9NJGlnqotywxy5cLkP3wB
Tq56lGN/vqiBWA7Q/u2EzguO/GX0tUELOIRuSyTewk7vonHGFG/Owl/lrP1ooMHO
WjqjF5JKIuen3gVpYXNapYvLUZJsrI33Ya8koQP+qI12ZlJfLiI9CngW+D/42RsY
dcg1dgwk9o8qMnDobKYOGt7uftbT6sS3mS+QTw6oGjcywxULVZyTiOtmxu1wCkQz
BkkNPMC4uQxChkIBzwOnEKpgs2GUVCsCYJ0FgMTwF2IfUOCNFZAj/uv4i0JDEhhD
S97OirgZZzFKcJtZJ1uIyL0JNp6cw2uESUHUjTR8iSTTziAtU6e2goagx9urG1fE
Glmc9vMIQBAlZdBMmwpr1G1qmLiZBnsEWkkQYmmr1CuU/K/i0a46TYN49DCAG1dh
GPRtV1zNact2kyldrQ+SzrtSzm6P1xt5HQV5Q2Dng7kCvMIFA11GfEMLjgx+DXPi
ty/p2ES/0f0s2Bk21NxzmJN6wnuXn5hsES4XJuthOcQtmBVYedPZD+cteF1WbeAH
qo5I25ONfjlEub3/yw0Yrm0fW9nwntLUQ7JQwTZ6kEBVpRIDZESaU1S6F1axEcaV
AiZBLD58c7DFLPEnZC6vvmzpgoHdczqU/hC9GXlf1mjQmzcr6oL/SV5NIbzqD+f3
GKcJGXf15yGCyJjH/fTt2SmTOusAbcV5RHFsyaeuJA3nN72l5/Jf5Djjf+loijUQ
q/y8NcN1ec8DoaD5BaeMlangdXcYUZFUxbBWkYpetVbEZolV1dXrqAwC/dVo1zxR
BKDAXc5P+6QnQLqXYISiJLXDR//4Q2icEmTR4Qea51cgqX19HRdh+JbiAsEbdrbR
1UWOA4fTFNS48oi/uxo/Fa/63NcF1rnuKRbdg/jq8GLwzKOusyTmltvhgZBKPQje
he50uYnq1/LvgpUcvintYnZlK8uvgTGKzPtK7EFF37Jdvzw26amVcCCds5KH/fR2
jBBpqw7r7C67d4PKQb8c6bN/RcLZXqrBd7dMvdIVZ2FhSYtcTOpi107WjwD7nQob
ptJw/If+aRC12KEyyiH2nP8QeJUiXfSvRKLQDr4J+6F+Y394FcA1uBWWFBW4bs0i
4e5ywmOW7+ImbMq5D/Q3WBDGGVHQnfaNByRacrw6OtWDlAQtQXzBGdcSZ/Zbr5We
4PezBpHczecYIEwXUrKSOOalIcS5OTH32Jvym1Hz2rPmpadZkDRSrWTF1a5sWskX
72uxN6K8153vJk4DiHObeSi5/EGO5LxdnT3Ow3+oZCbTDo0C/BNs4SIGr8rmwslB
8DK6j4CcUmTlLXCu0VnGKVlYWq7t1duNpei/HpERWnl4Ay4QSp1ZW9rRl7tVtHpP
U5hPy/U9s7VexP44NusKtdVqn/20meKT7ohEakS9veUqAE/CqYPqEZ94wi9SVgSA
8jat9h6iEhOvTFBwbNG6LsjF5Tlgfb7CFHOr0WZbo6IofHcvLTercPWfH0b79s5Y
dp7epN4rmsUMyJD6WbjjJmLWYUcHgifz5Yq1T0BSGoZ0IACWxNDaUVmLjzCrtUQ0
eb1TQkfdj9DBboWBmzyLoulbg10yaBd18lo2nq1250skQGZLASiDDSMyKfNGeO7u
b+HrY3NS7NLaWEJRa+J8+pk8XjcajLbKZCqFpf7t67KwV032ZTEnuU91a3sj44KU
BIhmRVP5vlIz5YVXa02jI+FkegW95RoIpjSnoMH+19K/j3x62Kcwwrxhl4SBlDoq
+ElFAFAl1q1ujvDUt+6F4L7P6V4fE12tMAN+tn22sDzeIgWKbjqf0cNWFY58ag1s
1e420I+edxIfCdtSLliL8vId7nEOiVHussvtDngdGMgYTx5odcZJtg7TLBDaMvu0
sBXoLszVk23HvGkghxI4nnRIdUMbgtRhnXFJfM+oFuqnJw/AGSGHimaf2Cwoh/Hp
MYFFCI/2aoMZShJffqD+eLyYBR97WsdeKK2wRXThhwxT1iAniOd7FjtD7b881dYE
8UFTXdochYD5zNDj69hSCMdcojtz69rBAMG/6lUqvANXvxx9640uzqZ18JcmsxtA
U2MCb14EUY01TXNjIdP7gIwFJrezaa0QuCcSmhoSfcVL77GUSAFumGD/+gOhxkqA
se1OKn34sozZY5F74ot0hkwZePZOB7luXkGFHa1qrx5NwQVPJ3f8tE5yk+67627j
eJJjvJ3dOv87/0HwjycJdN2Z8Yz2FyaW7sX6j28w93hQJ/4KokUJ860gokxVy5zF
Gi5j2EzUnHiYS0ZhNCg8yE76xzDCkim1pqEm7NSkL54KKiYVIDOiIqj/4R4pUp+i
S76JrolW/55/nhaQ/Vk2SAcpZHXVEJGJBKj2H6//S7ilGz9d13bB3rby0tjBxvMH
vRHbx+dbcgNWJ4EeWd9+VLi1j8HeOqcImqu/nMTK1Dc/TRgNDIqOQhJ3rR8Li/8l
uDCq5tEM925p7g2+btXJhkktrZcAVE28RzLFg/zlcC63QaJ3aihuXOZspoYmhUbg
Ii6rZe46yw++pRjxfnEPzq6Ekag6Sd8ISC1OFiPONuvjF5vWvVXDy9L1jFDw/9ng
PAmTBRFfL6xeTkH1+uXp8f+5HXM/p27RbyfSToyGtym2ypnZeUunb7HUiWRDAbld
hG644R3Tioi3nlLrxaB5klxOWUqGmCpa547YYwa3bzclzY0yLeX7M7gvkrQNoBMa
tDsZK/AYfS5nJ6/sN+wGGGrXyLI+bzEOPOC7IdGjlQs5DwYUtj4Ycu1ELQBIFXeC
AtiPQcflGMpnN9o5kzwb1nUyNcp6/5YCb68MTrK52743e6SycfpRaa84fUKacz89
UTt1ZqL5vgleWV2bEVj6BoKrmdAF4bAk6knz6DXKJ1Kes7RKIWFC2hjwlvoGuNlP
p9524uDYFbRNN1XYIK+Tp68fcha1wK/PIN6Jk5ul/WrmyjlNCxvks/SaKEeYiBDB
5Lmkb1U7rJxiEwdQEDcsCLHbOx9hG1ssxbGwT3la6uq2EaaG+9x7Rr75ZpA1WrZb
7S3/SzEjZ33s+iIzEWq9+RE9+B7DtbEeDRMTK1Xttg2x6rhQsa3kY3zAmV0eB01H
v1R1A3gozyz+FvaOU2j98DZFR00k83t1Onz+tA8QexcYQ/ZM4NYtsiuVfW9lYnlj
iGEaku63VmhRQ2p/zGVHnHuVTLxRudu7o2+ToD46KPx3njZL1vZbJh5kg3KmMOOR
874AqyP4QrrGO1r5Hw+RKOkdi7OAMZmLrGxyLOLDeQmkv4moOCP24x4FUmM7JqOv
1TIdU78DaIzhX80I2k9VrtRWY8k0Ao3JsJkozFIEtx0bunRBMlUkLug4ilGfySAJ
d8jkyZb8QZQVwv6KRR4phczZJLSnYapbt5Rojg1dptHyuT9zGJyUNapfzBrXogwC
LZi19eD8ilgV3NRar9X90priG1oMtEpPw1ZAG/3l1uV3N0mWe8yrPbbtmV63TqIM
WH8sBMBtSKetNY/cj2KaXirgqfALnLNuxuEjKvpm4bTJFN67FmUMZgaPnkGYGQuN
WTXHkKBv+MFfZh3MQryAGKi2ZEpW/U4H6dVF45bo2HvZMvt5cNr5VH6jxUrv3KIJ
CdfZwrVfB0GpeaFrudj1ej8sAyIDn29UrP891OB7VLf2uTMkv8NKWJ7QyCg4TwNa
vjHLPYhitwg8iD+jb2FL8TvRcaVnz4BFbJqAE1fCh0w1GoWrBwdFqeL+hOXg1jf/
5mRxPBrJDATdY127hrNY9e/439T9JoUxoSbyRdNeMktAgwung2sYw2d97YgoJp7E
wiRQdzBrR0/ZIpe2+xrbcIlz3olNQY6H2e4bofSnpXL4dmTf+lNR6J7Qak06BSO5
WZqvNjiSppr2jni2/UMccZZCdOgBKHp0v8Z2VWf9QVhSiYaN+MBZEg8mOQIgR+vV
EypxiSthNeQ4cD+fKsnesz0pf9BmbyFkLVVUJnsEJd8afu57rdU1U/m/Z6Ek58s6
4njKTr2/kWPwxfog5dS59D0nLntwT0SJa1y20j58gPE3kyGM+OiFqPPM74mdiuFV
I/2rKo/bj/e2TfY7z/8CFXMwHc404lxJwOYSqjk/r/cJxn/AoA2ZqRI2CHTW1MAz
zWYGtagv7mFy0wGqHdajbMRB0ShA7fB0gTZluqKpGAPH8inlo5R1io0kFF6rSv2a
J0n7mWQIYOk7PyC/Z3Ixi7LOoQQTpfCxpNTiXRwZh0KmfsCmZmcjOb8bQLj1yvmv
h5zXxkUrHmFzz9pab0LDThFVfqnPYoq02pG43YwSAjNM9m3MEI4joP9V7khZIL+1
vnM9zQKD2rHCGzUiewsw+GFV+4SYk0ZhzrRRrHHDsbKcMZI4Y0oj1/BV91wIFpIN
El3WKcDytw080uMFDjqYiaKtf5oGMufSUicj4ZLs6di/rdDqxFpZuk1oeSeJ/07J
QCOgo2pnDCeVt3cMyB0hxLUakSe6KymyIfXnNzJRxPChXyRc2d5E9JCECM+c2e58
x7SihTtX3qq0RcVLVmo5tFpaVwSzwrTCgBLQKLAO3MqrgM842GKfLqSomSoBp+C5
TcsOHr7IfLS1slCeXl0H1mSA5byYvy26medGD99g0tcsGR4R2VelBciIKDEwZH4u
ND7Miekv6sKL16bmOS21Uer8SrdjEDC7WKzUwBolScjW1FtZMAlztFcqm2T9vton
P3Gvw0WXqW+7NQAWiKNjcD0FxvoZ69cr5zYI9ZduGAL9dneWL3GD7ab9+cPzWE3L
XVueBBd+VKbb0p7jsvjx5+WSyu6phmvRoTDD4DX4Jx/KEu3ecwr7r23pgs/UTHyC
4c6jHqG0STUcgGCiPAHXRrRahFpx0o6FGDwQ0mSy1C9V//F8mY9u8CFZnJm3xJX/
cI2bJWBf6ua2Ac1nESZx6JMFJ5FBFgLjr+O5qAP+yL13l9Js+ICXPsiRxYpoFKxC
EgNBjiYj5a/MXySntmZAPoBeADfuHK9G7SqE2RQmVGrUiy2neloIz3BeomNC4ciZ
0E3u9SFOqYRv6eDKAOgBwZNOs1QzQJgzST8ro0qlzsD+lBdVWg2SMNybI8amrh22
Rgp5TxEvtLutfNWNhjLQMDLKUA2xPyNKDkXS4uHWpApCW2YZBTmz9jL+iqEqo5BX
7N9ujxAkj1o3WvrZsav3C03xNHBRtXaTnXF0K3GVzPQpmSn99Gx89DHmSobdLp7W
VjiFkHP3zSutXCIBKQPcnjoSZ3I7YGFpNzHeIFQ4JM+gAyDuqrO0yw5MJJMI8ulJ
KprX/EaaVgRLOiCyzJpVwQpidiqj2geK2QcW2JmIWettxvblfXFfW9g8feXxIOsh
9Ovzb8sPoqsdcZF99rpv038lTvK8hLRpIG9rioCQRclaWWG3DckNR27LyFrRBJ5e
8RqOfwPSer3CcmTxdKxW8E6Ccpu/Qah0EYbisD3fUuWYnKTUbpYFQAt+SRnqGkYn
TV/k6Vo+N5fXTr8SkN1iJ/+jz5ccQXAgdX9k+sBjrrmKmRzDPKg3V/51SRzbcnBD
rOBSMr9ioSIdDeh+Mu/haOOJXzZ4sQbmyRzr+AqTwuS2Wz4tj2WA1WJjSd6FW8+4
bhI0AT6T/wf1f8PNncZULs+SA37U8WQqbZUDkT4Y3fLoYdutxdJHM8OOOD7gbCrp
pmyU8QZ3YpwPuTxa3ega2JY0N1Ht+bhlUWq11gQkyGXncf9sGCnlQFbuikTI3Jk2
qhMC9N5FE0w8hEyf/L5+XTKlIx/Fv7PRcG3dzavqmRpO7VHjZ9K9IE35mUi9Psw+
8/F7r1jRpya7DTiTfZ5XXZo3RVAJuwFVxyvoD0qeDUM6ijbPjC6tXXaofGRpD4JR
dDN1p/QNuOeB5wptJWjRwbXg5Eeek7FHX5x4gxPWAXK6a2G/I9GeGZ4u0BJ0DKPv
++rrpm5V0W9pm5r//x0eJpNpTIfKWfM1Go7pOXncZOpBDGW5KQy5CgsT3knUSIHb
O8wCqmW1tIwuqHw5KEM5O+BSn3fydM3DKmvQ5380Xtr8KnEsYfhhglg/g7SXLf3O
BdRWCO+g5kCEEvZt1X3ZSnRWmKn4Uo0V0ldPZqWUQLMQ4Duje1ORSlTZKA3lH5DC
lI5zNwI3l7EOa+gdAA6faF2slVDYHvH0Oxns8vEwYzOWnYjBXz8l8wfxOJeqIZMO
dShtaO3t60XjJMFDU9+rwaRmKWfFoTJPMYcO21p9OkwMeSEym7wiPNq9zQG4S9ZL
nbU4hN3tzSG/0DiImPA8h41wrawHG96FwuYUX8vX6VOohhw4fH5MwWEp4gPrqnkF
LeztqBywTb/1SYTel/v0qUVOOMHNT0gJ7gtUkgyXY4SjCkX7oSHiQ+mSJLESi0Ny
kRsjtgIalEzh/6es4rIQIF8Z1OrTmPCG7MgbxJvSlNOoFBBBAFukFVmx2ciaLafu
KYrtGen+H6/n2kMyS5C5xTBzc2ssjT+BnXIubCjYNOcrr3/wanvkGyXoHB6UCvQi
9ExbpSrKwjVG14tp63FJKMoeHD953y+iziVG/X8g/gsVmnZBZBN7g7kZI4uXRIP2
7sR8W/kyr6YrMib+ivsyJ9ZjficNj04zTZaHOHankbpiO5Aor+BXKCnt3EqbctkN
Aj1437rZwYMX6B1Iv7ENn9qsGFRXALflVXgOspIT1Y5lts7+Uoi5WILPG0vn9Egq
HtciDXJK2KWU49/yFbtz87yODejGlt3i4jFU5gysDSxe25hMI2K8gX5r1i9YwjOw
RJQkSsDINK9tgyYpf6KUxjbKKuP8eWnK21UVZGsFT4PExaiMV58eb6uyExDEx1cM
S08UgZ6MAMij+a3TWntHcdBY7dB15oTtVYPImKIOW7BOPIwpRA2ZPl9sqt8BlK4G
5e94iPBCy7cfjMgyoU4q5a42cb2+Q8FbXL7nowu6tOa9BJ/lI3nsVzqw0R0axrOO
t370qdD131PvSPGF/cGnzOME2ov/4w6ZHMnLYcc2aiv7b8EqmAtziWQ/OykZf7hu
YDAc2BjzV6mO5Qjw6kvnnkjTVgrm4oKl3bcx3E3ni156Doufiv5x+qBJWarOMvep
vU8/L/gY3swfi5X8zF5yr5kPVbC3N/rrVPrxb3vVqa5wRNWq7CNM6ZitQJ9Os4fe
4uAat4eSt37bsLZV0cvZQHAHwSykWXtw/yk1UqiicjZ0YE4tFy5rDQ2ZxMfH+htZ
dwfYYdlYGfHGntkc4QPzrttCJ5AMLyWbicIW1csv4eOTfn/iknypdf0rz9Ai3eIf
eo/x/2l5b+myAp+RsgW0VO8DdnktUp/E2YxBgMb5s9YYkiDvsG0QsgR+EiV03o7I
TZ4jSAqxUj+90ZEZ6M+i5E6gT8xi9LqNZxB8HH4uPPXrtMZmcw9oqa+fCStONqBj
byxkpNFYR3MAeVYnbd+8VKrAikAsMxvTRK+uU9pQbBBWWWkX9YItUHyCBzopkP6J
OSGi9EYjtU5eeXQdhlMVnOfsB/tGgUlZ8DG5B/TcbqFaSRVLAy3BVtjat09r8rvb
uMfgk756L9VTQyQlwaGWjX2Kvg7sbkhr/dY+DD7nQIbdYy9R2LUTfUH7FBd59TEy
OSHiz8HgNmqOY1JsMx+tI86GVVMpLe2VVDjxDKD6EbFcyN/f+Ku4MsaQAh6HeXPP
Q7h3ZVjIpcnJLbnQ5vI7yX8gllzITPKnN+JSoCTJ+rYHhKmqnNmdBpmPFte/WaHK
BY1X+TAaGwAUKG00/6A/IvGbEvjX8vcyYlQWz3NO3yCBTTiQybbjeOW40mjTe9Q3
267oMAi/TJ7g3eEZtloGgrh5zqAyc3BrEK0gEyrN6kPT0a2MRrknvgOruM5ZlNvG
4g4OOz/rsRla10dxAWkiYI7Q7svHHdPixz6Z1Zpg1Jhg5YaeC60155SQ0i/Y7Wnv
qxgPuyjFDI9i0Fv9mU2MeOdgWurHRbHa5QkIkfxest2mcrAueuPOLc5PBrOZEnNC
jiNNnfL8El8OzJXNxUJUogluyEMZI+AFHZDsnUB+WIWf0RppBCOVnB5QxMXF6vXE
0APPZ2BQnpWpyYwoMgru7tBg02fPccEr9AE9Pbc8wJYlZSIO219sIJzbRtpL9hGj
8bapjeFSiMyUZKPHRhpeEtixTFLrHnbwgXU6rXkcyx+vzMwMQoVNYVYjibqsALBo
lXzrWRpU8o8QmKxoFoThWNkd0xhVY7XOJB9gFNR+B+MCV8L+Fh4da/pks4ALEu+P
/Q4w+D57skL8oP7HcNKTAZosBphESU5hKDDgJxCjMgzCTOK6EvDwmJkjgNhMe6LX
75ueCc2aeJI8Sf8RS858GNkwjoMWSuJUZ+v/yjrH4eRX1sS/ZObqKY24Qip4GoxX
Ax52INP/zAbQxpDVXRfk27tYN1SesJmotcCq8wdngrRe0998ndgws5UxTUkAMMbH
Heh/7iTY6XD01ZP0J0OEaTGTDg/vGJbGw42ik7NJTeI1zFz924YI7xI/Cy4K7cL5
GRKEnomwQ7BsXAlp7FvT1AYw/3Bn+1hGuPSLlsdN1YYuyEpsXtGSun5siZl/X+R5
xs615NTq+/a7EgoJ7ODBwzAdKOkYpMibG6qhIpdOrBo3cstMlsUs7DutI0zsyRoU
oj5kNDQKqZZa0TBaDuOwL/8SPzcfyETTLly5kXMqPAAUxdZ9TFEMmqoVVUrcFNO6
HXDeJudgtIEaurtWzWM6m4znVuEG4BngjXiKh13c+ev05yiDOhyItEK6m2Um68Q/
HNVnQrC48UQcOM+DCnwX9YpjQid6YVJgPg5SHLHf47baz80vYB9j+Metjj3jRRx6
uUJSNIX96IYxI1971hPFsBHsquQCCSQOywmIHbag2tvPslh6scz6hU1MlyyiRbL+
8WfiigwLU9jDu14qlO6b5yFYvfTaUqlE6I3qFNXRnH+oronGBdpjcOe/sM781jzk
DAnJFhNhX5GBMVqWkm8fCRnaaIMvN9XNUukZJBqxU5vnxk40LDTyvDfuuQIXSE4x
FMnOn8WxS58g1xzFnrNScNCcwPFQf2Tey0RzyB1E+Q7act5NGHtxhpwzl9UX9V5L
nnOVo6rQwLoFiB6nBEp2+9ror3OvAkUQqvGVAtxXk/oFS9wQ7FTTExPt7GqrM6dg
FHSRa7EoFWIMwmt9YXjDWkkbEcysksGS9gBITxXbsVxTHXX2c8LNnfrmezEKliQU
qbWr0opR87cv1JS0UK8aWJdAItqfNkw1cfqkLFSKos4WnizvPwclhVcwgxURd83t
l71Rwlj9acD0xDpTZVeNhTGRxBHastOimQ/eAgKgNA+e+Oqh8fTderlnmFdV+y0J
vl/9B2H/K9ugye1ExjnQF7OnD2bKHIjkz4dbRRISvxbMbNLSVzVToF3MzI6uVM+t
+bS6pq5u5ZiPs6tb/ODLtrijJcZcn5Zfp/cM4m/wtvIO7/U5PI250nIZsIQ/o7JZ
0DVZTKJkdyCarGdX1d+5XSFfI4i5z5x8OUrXXb7xddb8Fg+Wu5xiRuEPWm95EjaX
IVf5IqJRLYIhshJ0eweFrZBd/de3IzKh10ZNjcpevoBf76PcwUUXpqVgDvxHInjg
RXtT53DO/cxLBP8l3RCg8cWKHiqFbCjdpNCb73hJfJGdC05lSvoFg2Kqs/A9TM5B
WzAFTQHewG9Z+xhSjAtb9L9flJlJwajl4hQWDlXODmwZ1UIbG8c7W44WNHcZYaES
BSfDYUNx94SqAR51JxZLg+MuWrM6AB2ydm8a5ucBhxwlJxa5s8L53yuRPfH17xUm
Aa33h0yhDuoZLYjSwBSw0MyLpFCCthoxvKz4s39DL5y7gUx0NQ58clqxvH4VVh4N
04bk9cpiv8PcdeDRdgNzbpBMCmo1i27gTdxgKdT7D7hC3G42YZgaTJVT0yVvMw3q
lVaw6zX58pTNkHCvuSvveC++v1Mniz4OwfD8yrRnbNrAVrqBrnADfcWvgvyW6tkz
RaP5YYwimTIYkvzw3xS3gxyhY1g2bdgQ/cybtY39DTWx0EINpDDj2BD9+C+ToJIc
R1XwORWa5d1A/qWB6CugFzSvhmnyomo/hESzyS37CoU14RlZTXbJrp8kyRSG+GHc
lQn5s51I+4LE0YzI9VvVo2XeXx++gIt82bc8VYz4vUGWhMNT762IkJC5vKT+A5b9
Kt6OZ9geu8EA1/78dNl+arjOW916cyjda45EdOxpaV8GemcoaoPb2IkFjcMmg8bb
dIlr0s6CMzzjk+4rmOiKAO20zjHg+LafSEYbhkxPlNqOYEc9+F2P9lqd/qHALXw5
z2dEswU0HBKca7WWtNdj/eGJdHy4O+kMDvAg84hTCqLcMpQGhcUPtO5fUl5PZ7a8
eAUh/KGARf2dRu32+7s5PJEuMjTn9lX1OqhX/1Bx47ni1O47cg6rer9W/mLJbSbN
NqU6lQLJ6qbJTO10kcep++8hcV0CTi6zDhn1M/4xsgeOXIhN7aARa6/WBPSNxzDw
h+T4vjLY7hPWTkrX+XJqUKopI3oqR0x4GjrECVYjNoAyMLuVw6aytHPBJPdDRGTR
zqmOn5CIwfPklOa1B1fzXqq5dUmyaEkVE4EXQ4/PIRc5ttcnS3zqp6NELwD48jGY
6B52zYzBQgycuWgcJsuPsh0TjWHPOiG+6Li9vcAZ8nwVgLex7P2yI5ANUqwakwY7
DHFfRb1cfSNE4RlCT+B4yssKbmn+JleVH5LBTmSbm4LBIN0Vryo4XK876DPcihie
e9fi/MeElnHm8d1NiMtD78Gsbaxo9i8vlYDKHMUD1cfQxCxc7oAyIWL//G6Z+ZwX
wweP+zDfYc+lFsXA85vtbxl9it/wfmZUoWByaBH6lBd3oBvuGCNnTbnvSFPhkLZk
jQ789jzroT+/qGGibWSvLz+d4r3X4Jm/kkL/XKtBbBFg5E8znw3nFQHAmDsijgyd
eDZZ0+nwmMKHNdQfRcnDprDuOgXI7IVoWj+jLVeh/XpCmjk5nyPD4IdqSWXnka8X
BietCdxI3E1dIyz2RZOcyhrDOZr7e07Na+xW6tEO2rgFmU+AbmyIUEh1VoyKYfb5
LMSlQ/+47l3CctFm68D3QLzTAZrUF4UHSWqEyiDcfkEgMt1+NHgQBiosy6fATAYw
hsrG5aAtUb/Y9Q4VBNewlEH2WU0jTGEas+2z+NJcG3pnmgiC3rgKtevJc2b6ygwS
tzMH2MNIGvnkCkeJ642oKVzKUiWUit4C/VHpxGPYesVbAKBlSWTop4neHfEACH9v
/5Js4LbiEKfgT8ZLetikZQ9nvbmKA50MLuLiaJdtExu8daZCSNWQv4Rw2WRdlgKw
MUr0RT64741ee2RuzdPov8+o6m1nV2MlIaNADB3zXp6rzmuxcoBrTClUMMlRXDMC
Dn9oQbc2K92Cudv+8sMMD6E9yKGgwqv8bZDRoKJ/r2nHGIFHuU3fcs+CUdYudzPD
V8x+wdDbA3QisJIxgw0BVDxT8BLfF3/ir2Z7NyxCoJpcku6eQvSBpdGwz0e7KTcF
DHOcFUBZ+MjfXb3fHgFozYrWZ+9HrAZxvv/m6aV/6AhgtZwOYIpPXfJdn/LqPvjN
OQeoxyeUZkw/nJNeNYl7BwseuZyOD5L2B4rbUFMlu8+fflJLdKW0bVsjWaOkrZSh
da9r/Mp5JG+4fWyqE2Iu91B/CSqfxNuLZYQjgHxgZua+K7fUf73ZSj9Vniwxq+Y6
KnrlrphNiusCSUY+uuBjmBk9lIKMHw1RcJAcIWKXWBgTVVCppTzFTM5G2TUo/9jB
eaTdOoellIoJvsErZUrPUqQdDeXUNJli+3Vg6B/Cpi3PI2JRyh01u4mK6Yqcxyc9
y5JW96bHR7ENa+UMSHzSzwESxQKLn9lsRta97DNnya+RFEjQHXqAQYK0fhgKW5VI
Qpy4nHPo0aabg97Ei5Nn2uQQoQ25FqbiQYbUdnmSRgEM68YXEo5HSJ8BSwqPWOdX
c2XDpLdOIBOk9shpSgIg52ZmZJOQK2h3NXcIfU7TG+GwIpG9iPuDQ/IO+2eQx2/0
vEyPFU4kvroaAA2L2xIGHfbjvMXfdwT70fwYEWZUSHDpot+I0wUahKl2ZjS7VHmn
pGmuSErKO7P+RW78uF2gOy5ien5PuV1j/4WRhHScdmRoKPf7PBH5D1kaNMvMr9qd
vauspolbTTlNpKwAfkoEB/QC56U8gD8tz8ZW3G9DkQEJj5FE1q3+WLVzBS2dl/x0
ECMzVni98QIKo8XbgEvi2SWsCCxSLQ8TrZSUDQg5OCdo1xlHxMALC8fFH6USBdIn
Tpo7SjIREJ0yk09rO46OMEr4rE2x2DuJNNVnBESL22yecu3RkbaoxleWB2PK/SA/
0cc0DYpqHxh8GUSB5FcVeWGFlM4bl+hDVS4saklePrkIGrLV7dTR6Jvaw00CuDWO
r24uLqaH5KTTA5HG2HH+02wujkJJBkLTSjPzhaHT76I4BwaOllaK7az25HN1tC19
ZIH0Gq3KfczUHyD2LYBLc9SXlyrURrpwhClc6yzih9TE5FtIJnI9TIXt6kuvC5Is
a7DnGCVZWUH2Lq4dpAEXT36EhSjWCOnSKSUYrF+zqzamaCEu6+QHrV8CUvNLGqCA
VyAf+seQs1az++SwA0dv4zor6Ja2+pFSxdYP0ljphE7Nwb6YEhgDybFqKVoWphMY
MzqqEvl/3WwOGud4p6tS7PQyikzdD6CqQpi6eIAHJYVuxBx8GXQFkduKfGfM7F8B
bVObCUOMM9teqWQWCLwttkp5qx1pxNjZOc6LeyJHr4rX3z0o661m7wb7XYUdnGZG
EUZyMl/8Q1Iv4e43he8C71Y6W+tS71U6sSagVy5gl22i8Z6dQOCCfbpmMQH3Boea
7DI7n027gDFzge5epz4Ys0+4NaZdfRCBTS66KZ5kmxopMjFOR3nMdxSHrRRZoeSL
ydkvYzQz6llBwViUjOUGKDfpY1xb68leCoxCvNqObRmx/X8TugMe80rpJyY7Rzej
hFZg88KdwlxQ+DL9wYvsuwcqi0kK4Hlc3khkXk09zkWZKfFoIo76kNjrIac/HHOP
iK6PohWLaq/fft62HXOpHSn5+BvLkjsSUbSrnKNmoGDISopj4nvBZ3NJ3WpT9zkD
Vw/2zXiczwcdpbrIIKep5I0J/d2QBYVsfCiV2bYKaa6VOhymZhGGCRNJAy8iXpI2
I53Kmwrb5OgTQrjxNldo4yzdCUR+MjQ0VzzCKaaQYmhVux5l9Ax+93HLLAfUJeQj
vyRODpSErIKXvT6LAPfRsIBy1Hc7jgKg6abJcazfR8EVr/MkWqEkYkV2tbMhgCd7
FQfWIXIvnoXH0daoRPG/I+h8BcC6wZwT3tQnNppclLhC6ky+A6Q1CFCbsyiPV6Hv
Zn0I6dbjNGy0w4zeG6cqWzgBQwk9HPfTe56HKJ9VGnG9K+750E/aH5PWtkllaH/N
3ruX6V4/qUr0HWtPWtB0GiTuLX5SayogTjKbBb4A3IJ1bIinyrZidXkuK238bn6K
Sch2UgFv7BZqEF8xGd5o829QJas0FympkqpPnTw/AlnCd9VDTSpEzueVtqYXLrrX
cl1ht7Wp7nbK7HzcizXW1+vYyvS+I56qDwjBePButBIijmCPqKPUCn/1Ody7lVUY
Fjl71lof/iEynfJitASg3PrYKef5VGrcEKHJnNtNn4Fbtdip9bVTe8cFk3LcEF9+
hqs3PZcW/GJRAtLMUbVeuucuUy82cooDNS0dpR+/lVXwSiujrKxzkWxDRO0HMjZM
qpUvLh1vG6DwguS7KgW3Y+oq2+DzBSmzQCJJWqtqZ2Dhw3GDLtZTWQFnrjnB2FCH
zYxTQrtGlOmQeyQVKAFMHqu9DUMSj+Aq9fhpKIzwBH3XoAFgflmhO1XVcAJXqQVy
Qna5DLmUIdF39m8gLgfWzpfTaHpPYYT2P+h4eXFsIMClq7C8rmGyRRPmB6RWIUeH
xmX1eDLLqWyUnx+07Hn33u5P7MtO0TDgNbBVnovW607sTsh36nLc456vNFsexRfH
0cjYe/in5pK4gZNSguSaxiS2CHCuJ9fGfyqcS0Cqd4RVewjp1hQ8LgXBINQAAgVK
6P4gLWDNF/QGGRYUzSniumRIZkglch84VApCDx6tblrxgiZD/ciQ81f0CalzjRlk
QfdA2zK0f79vR/DwlQCIM1ukKgKgkCbQXlJA3DSqH0/jcpnRRQ127G2EDIIkO4Zq
aVAgTVOlwTZvOgEBMfJwWEnawXu6w/a1IiEKRK1LgDhWiVrDpYTHZMUEBvYeGj0C
M4wO9qMKf33tbRjUtYHR6/ei+4kNyAoyeEOhrP8Nlf7s+bhkcLQMfOwRGwUUntgh
5VDc4/9wAg7tJl5M1OET4QIP7Ec8dGrCK7S0jO/m6wKqLBrbKm+dt3vIl4A/r0Jc
Ft1yJJkXIM3wI7CyV6BxV+rpJ3//K27wn5soTZutVDAH8ZoCy8tbwe+uRwDOeEeK
mIXv32OrHAAAof3EN8+cczeLI0h8PCfl1TGoBxdeUkyd5yGO2TvwoNKg0tjk9eJP
kB+0qhQx3vILrOel24xeD/ScxmonXcdTvlHRbnVwPk+8Kj/HBH9JM65INRU3MWsz
IpwK+Rxr3L5xvoxyOoWhSa3Doz/C5uFrkkfByGmD1aUML6uc+IgsJusJRF0TICxe
njtmS4fYD0aJuqDAzI/rNbYlcqNqtesSD0hcq2jB1EBJxc3b6CyrfUmfJ2fTQdLO
atwYnmKmI2zw2/BoS8EgLHw9d4EDQ5tdsF8DhyR39O5XD4GgRJWJ9mBzH2xz7+AO
T2uM4ZSiYchxgcKvBOUi1RAf9kbJ5mk1vADqwExZzhnaJau8mIWbe7kVYrsvshl7
r5hcs8ClZohsDUgsFliBjcdrFR/+wPfumPd0yxQhRl2GTMipgRvvbNyfMLLPZi1D
aGSiQF5q0FyY8GlCOIZAbDUmeP6rApYr9JrNaFCBQXtIY7RJbxskdPHWGjZxNnB6
iQj38awOtpg5CYQC+2PcyOas8a7PIwJfxfv93jW8Ap09r4eoZaO2cs6wC79y1oa8
HJNZAwJFAlHrYDQOEdHbw03ZkGu8YGiV/AwLIQGRVirPp5/Udlu1RqQHTsQjbavw
58d4eKWj1Gy+nUpQ/wnqxcH8Kb0gLUPkcv1ykXjwmZEqFm3XsYAfYfmwzzH2mrTb
Z0eiYzHoJCLg6GqTfWByc5oCS7/gfSf2VLO7FrGVQ1Kj9QoIRNjGkKiMhUPTMeUt
yciE+fl+IvMoCZHNU8ht3AGhea6jOd+8Cc4JT7blrPZX3gIkUgLNHyhQMCVMyBzy
s2ef/OyPo0k5PkZZbrkeB2oiuSvE+FWx6e7teS4WxF6yAyV5/EypBgtNdgiFG1SE
/b0f0BP/ApqS/pynERjla84lXuidSmVg55bDbU+/hzDDUrhmhNwO/mnKnz2GROUe
/uCjRo5lpXDl8tT3DswsI1pO02EMD9EgrHUYnKCwbJOFprb+W3jX933Z1pel0a4h
z0NBjwQ8COLRjJbbV/vtDn6r7zb0+TKD73wcbXFaQtxK+CNZsu2IzZ4ukDS/EFF5
ceLvvqe+VPW0zJHxsCL/BiofSgA24seUiAQug5q46p8AwVzx6aVqWj/6B/mKuR/r
O1L+xRiZ6c1hsUfVSSkQ5X0V2zSzyBGfgjizPmRPJBaJL/zdW0vnvKN7IKGKsdVk
1YChq4+3fVg5YAwuZxlobGBpyQnLBWVG/hqnJEO01m3c0Tfpufg21unAI3HQ4Vkf
x/QmqaAO8EPuGnbdXXzx3LgFemJO7FO5bZ8xyzCMA2RUE1HSmmiqz60spdax/AZs
pWHE2CKxMy5xjQ+YQd90yRMQiuTX09Pe86zdrWy9e95zmmp/cPqxkENh+iabZVeh
Hztz755iEPXj8Qwi7ikrdMT41ZkuT78ESwIecah+oFxBsw16bikgg6b/dNol0u/g
Ap1yn8yRARKtRbsdugcq/RE75qfokBA3mCtkHJAzUFlHnqBAcxDPFk51I4fYvKTc
eVZAvHUG9aBAJFjFaMVRHqGIi2V3a9vwm+IFFp0daYmqeXSlG7w1bVDyy/ueYNb9
BE4uQ+jMvFzpmv2aiEQkXFF/N8BQiPv2eeZE9/5jpfueIHLLZ0p1wSx6X0TdXyF0
tIyIT2Q2ouAmztOcYgqcUCe7tFGS3HCbTTQjgpb0+7LjLeIIInDJdZ0GNG6e4akY
lTYvCfgUk4cVkStHsj1Ip1pkNzhycyuM6JyeDS90FdwuTmEMAgSq8BZPRZZFLY80
/wwngavsKxc1veWijMLU4IvTOvx6FHScHnWc5MsqKcxIh64cAxNMlye1IHWv9fKk
q7hxHgQJXW9DiyedOZLlP82s/A6oq6yi8FvFH9ExSBiIrlwbIOQjhRKtMKlRvVLd
v6+HhVzS3jkbUxILyUYxpGhPLsygrShZBjWksPl5b9+5X88F8NhV7JEYcTFOISPz
urOO9/5e9X7cDQLOB72gwq3DMcGy/La0gK57EBUUL8Cj+mceFxQeKPJfjzoaZvJw
i4exPso9t2WacyEoz8Vqq2Bn+ndzy8LZ+e+HnYHcg2uqtqHzZSbxWxoV28eX0brr
1fuPCU/K8nBZkpPblV/kyKl7aQZNtbFprxN5NswW1gcMWRM7zUYdQCgzjb24WgAo
R9oVrV79ekrlfAuNAC7j4JGG7gcIvf1tctbG9n8zRov7ng84Wb6oi0dtKMXHy8rO
43iXXGWT/oSqLgJbLGUNmB7r6R6I9uiWWwhOWOZ/pdZ3MOsQO3Y8U+jOAD6ZHMn2
JV+EDjpnL4Hcx/Aej+KkIMqSLwok247vS9g5+s6d/LfgrlBvHIgbv7LVXQIqmH3Q
dJwZ4HLf0BmlB3x4oMdoActd6AAsaRmPfu/wdlvuThPXCZ1m//JRR2VGuqyxP7c+
EY6rM/8E6xGn0Gi8segztR5osDLjQQEbWHZN/ELOGY9tTyUKOVl3GL+xR3eCiQhL
AceeVJA/84fTHwhRJap8TXfQylGunFMMH2rgvLpahhwQIRuWdDQ/BXlEzVpxKTh5
GGgYsCl/KSol/javT6/gATJTcZoHFqgRQXve702eaSkxCoC/F/VXEOOAy41uuobz
trF0XXl+dSmWBfyVS7T8p1MaQbQP4sIqG/Et99+U2ZXInLA0dpe499VAAUMjL+5H
2rsgGwlnbinPtMViqhUgNQCcx/aASeOOVs+0DX0yXZOmG5pK2tZUiO73C6rFzfjk
5cUnNc/1hD8g2XTcRG0zwxcgTL6kA92UlIDKsHuM53QGcJtFZAV3SQQdlziAVqvb
BXTXuCPK8U8gElm9V1LMib+2wPiXMDwUiZqIeG9H//dTjixK2NpHkTbJwLAqAQdJ
eyfIxgdzNAhfQHGQrIuZsW/LeOBuMSf8WTmJaNKYoE6GP6MoJNYTR+T67kCGafgK
AjXKlts4iFFPaTYb5SUBlbLBSgh+JMEK/TXhd1aPuV/imjrN4TKa84pG9oEm+A7N
/nT/x0sk2KY2DfKkkFJhD6+/+oWmdCUBChTBqtaNRCBee1aGIs5vMyXfBOQOpD0h
IqhpJsr9u6LqNgbHqxnhmg5iLab72IgVETVM21fgRXfjtlB1s+7pIE/ftePhkSD+
JTWuknkVlQt84fupf2EIpFCfbAwg07dqQ9lapUlg0049BFBJSUF/x1ctqNc31y+K
W8eagd4CsMBxG2LsmL+nDI1XjekF8UFbrJZfEabntzaLeNPWECfJvZ0y2sW6Bld8
nfxxpN86DcnZkjwkTiZmTiquv2dn5tLtqoDmhO67+GS1M4oX//GXcmiHm2vrVd9S
i1PexahbJdMn2SvpFTkRcOC8Y5tlr2qlRboMtu+0mbrA4nTFTxchvhPAvyMKwx6v
Pb9Pv5zRV/gGR6Cswewlds1Gx13pSjA/CRgS0kzvC4YR7VzMBqcJJhtqPrVhh8sd
pfLC+kNVFM5AyustR8NjM9ueIzEHRk4LYZ9O0/7fztR3ofjBrL4DS2Bt+HUpbWOQ
jZqXj8oCRZM1P2h4mXwBM0cMjdONPVEscdxn9vz45MEWJlbJp1D83Vsanj1Pt5wq
qKCssY/tws8SVuS9zCNQWu397oLCe4Coq5Bktd+ozv0xlUNjuzaTxa/kZfzyN9zR
OSwqKg3//lKPksYBh1nDnRGRKxGX4ABlLyCV9nS1/ToL6FeiuxM2bAQCgbV74fTo
z3q2QCaF50EwcqmOJrB+wUcy4pERadkHWf/FxOLAQvCGicdX7WXYSWN4EoHU+M7l
oHBScY7B2E6k7BG89q+HGOnhR37zR7nR4MxJNH4A1J4cC1AsIe2zzgVjw/P2f3P5
Im/reOrB/EA0wETJbwpsS1wfFBKcPO/8ZWH4Q2sCNOPjnN8CXgC6dQ6xZIX89Dbs
ysGrdYbVrIsVKbQEsoRpz4yFtklyDEzHxTxuQKzkwMHPT96ZeT1jSHUa7u7O/ox+
gtBt9L/vk5ifTORPjAxpzh3McV979xetmRTHubC9Gja6eKOrMLe4Fk+nTakcLiqf
n+JC7qKZb3AKlw0F0EAi+vA7VyvRB3sLEr1+VsVg2LOYCMgeqsQwia5EeD7nEiEW
g4KQeK41QS2ZDcQNqvJ5pWYVeTJ3HY/Spc/8i11qDOKwWNRRI06i0vC0LuDr7S1E
giFEWrjUwtYcn9A+sgERPt3v2wzBOe78Hm2RYfSpV+sdhQb1XZZnjF4dygChjbTz
WGj/J4DEpv48JywuEngy7Rk99BGw8lBkWRftEmXDMLE+M+bXVBODwWK0Yrb6/t5e
YO2qgVM1LUYCHSbR4dMPnURgikdzbSUZa56JmIdQk92HWBqo6TUvTzhKitPaZlTM
u5Aew1oQTUFQs4nYMBjshoP5mrzsUK17Mh/EasOtwCu4tb4kIStkPDVWT/Hu08oE
UXmUGFl0MAmxImYAQeSQZJndfRYjGnfAWANrHp+m+Ia4FRHiur4WOo3uaCMyreKt
Tqciy0eqaSS5+FlGCy9kBkeD+k+g4IomRm+iqdQuJ9Rm8IaSxvkxG9eABONaAZB6
l10FM5ea5ZkvXeIILLajFXble0UVHTWrGIocTz1keyh/cqZN22IC8vaENDsJayqZ
QDV49u9BjZSmc+BssUeKV/qHyHwjUVRyK8NO2NQ48P4Rj9z4w/syPTn1SwFjTGHR
93oT/jLSs+kV7h1tnxHc4f1VkiKaDV3Z5xIAz4Rwa2UVtPnmxsmkWdvoVReoZKa4
NFpXmqCkEPxTVcvBZFJ+0lwW6eXjt49LweLQ/tVgVTsDmF4g3SsD/OIBnZQQij4b
p9yQrgUbo3V7vvktDGFtjAOsl2Uc7tvT1dh/KQ/W8MZkcAAhEPyIvOgPno2LbJPg
MH2pFAXAYuolivOb/F5vkATNTpfCYc5KowQFaG0EOzpye2jKCQL4BhYE/suU7Vmq
56ZUGcPdcfXqelW9ofixFp90VKUXP1Zdd8by2fkwDJstHjclRCM67/Mf71aD2kRU
7wooo/sFzL/0CzRxQAFNy8YNbvP0tjV4GMoeUS7f1DgimEnsKmUY822E1VbKArk7
gzCxFya3Xkl4BsZBXXIv/6XpsuOaIX7d5CBSirRFXcDboqGBmr9SI3OXdXoWAoN8
ciJzSx0oXJOf4hudSYELP2JQzd75YEDQYciEYWss+f9LhN7T5DezYBBnIUWDrmdv
kZE+lLgcgzO627NmZa3lOsiigGJOMahlCRZH6tga8fkgGfB2K1vJvQs6dAUk+lKy
lyDhJrYw7hHh7sx9dWDaMa6YgReRg3/yzoDJ3BFtwUDDnepX+wxCKIIxo+zCGEId
dLysrSALBPuWQ/Uusn7uHtjS/TXnX5MdYsyP0ARV3MK0ySe1N8nLUM94TsdnKEUw
/4ALkueUb5Ep72PrNthsSs+C6TJqUiRTfaSKytfHgE6zSMhc03oJpzMPJB5dXfI3
CrHwv+BfCi5/V3TMtH02bmKvtL8URMPFE3Qvt5mbizjz7k4H/P8cASIRC7r4noIl
2D8EXub0BAJaV0Put0IWy3hUBQLUD1GTkGKsQRmVwIVCrMtQbVZ4TeWebKmJC6lH
N9+ZR8smXwJuSgu/OhxqIszBg2ASTTs6qlrcs/kYxPwcogwUxB2rJQBEATURzKuc
piG+UOQwOMy4LO0oYfEincvyhngocxxrvf+6XpFeol9HUNHflRFvLKulMRogKy7d
UjyOMyDQEGlroQj/xYlo2glziLVP6LJXrmXMhL2BdMEX6oveA5/JpudlFIhs1hAr
yW5mC1QQRDInSXT6KKqHN2HODn6e0b/3Cinzz7XmDs58pVJK6CaKViEGgJ6cDjm+
x78r/i3nPoo+RZggOolvVuWaFoTEkvUGgVXwshhKzE14Q4S7b1QUBtUteqI9GTgV
Vp146hneGWgEbW3be0V9YGrT5y6X9R0pKnxu83iNopcdRwdkRC7i+qsDPL4HVC1X
Mwys3PjvPZJFvQo1M17D3aJcSOc5gMvudS98OAHiUBPIFF5wMc+4ibctbigD2BAj
vfMtEnt9kyFNrgRJMkjJdIEWBl1Ofq0P0uFK4TDMHtn3mzafRqHJvR0TgylZf4Os
52ZQoD0/BAhEHqv052AyWd8jvGlr9RY5oTIslM+nJSkNxO22Hqrp+X+2b/R8KeTX
N8bpiv3L2CwiQr32ObRL9NhIgrEJKonysXe7NEgek12wBdwWfgD0j68Ktgyf28+x
5YjygwTjT3R2J1GNTv/BC9JL33sd2pLK8S8QUZAdXmaLGvJ44i+9gTykgVhpdrwO
7CoD7y6oAo+GQJQ4Kw0ZdcnwZ63eu/KjgCKL7/OTAyr5/uGW4SjEH90X7W4n8sAY
xeH4xv9KN4y1W6FsftHXefsyvcT3YUNUUNW+pFzDYxArnZuT42aGfWtXLJxyHDLo
86KhmeAmVsnqsA9iL2U4lEiz3gn39hGOr0ON8LD55NXPQ83R4UoedP/VgPz33lcd
Uu0Ho5yWxlK2Gcta9xWjIclUjXUps5Uy68/mz/4QMMXO68laqBvQ/hoDYfdQ8KLy
r8MB8RjCv9XCFYNPFdEXlFZmMu1JczUKTDi55IV+fCRkIxUUboLbEhe/7Mgt4p7f
4DG926HQet26A7csWaI/xYFm3GHnhZM61t9lbmITzaGADoo1DyexcDiTGBjmbcSy
LEEUnj+zlcpoBMhmdRCSHwlQ9WdDh9mVdiquUYGKumNB6dIekCZMZ4MQRJ6PKAQn
ELyyT0mftds3udCrHMEStI2SjrYlGtaphB1RjCYnaruTW7w/vNsEetFgKM3eH1U3
td3Mq+KU/qlvWWO2CvRdnFzvTCF8yjxU4dLCj/qx3kWjBa4u8n2NAYynPieIylw6
Tp5vyFKmE1fRLBNumQKAOxAE++m3QIpfKnFX+8pKoj/G5eBslYegsMN2hldzSgVZ
yzRHtDGRhAcJz8TbJCoKWlOFzNLLcOhjWcC5az3yo9UKdOr5jPc8tD3QE1nr+7Gk
Vw7iDMd0o+cq1q9za1EHpb6+I+Xp2DMv5P9wHcI2bpH0Lp41XbZzfV+fmQ5nNwlg
WRI/XJ8Jxz6X9cK+UiW+x1izRGFzfjw2HlqIta65VKfSYhy+xpUxDkpVrGU67VNG
B6DDzgNUtgteGAYQw7zb+LtCpKga8IZFjv7idmRAOWlSVsvCfpQdF4dGZ4/H9g1v
yTwX4NcK0PBJgbDFFq5kr8IWWTeSzPKXX7EMqNK5MY0SbZG77WC9xtNYav4hZbiE
ebu8BUI1kvCAaOZFAuS36yJ4/9aV+/JXjYx4O1JR17PbbPfXYiafN+Xj3wN32UeN
NY8nFLnla8UP4CFLvQiD3bUxsNZUtPCNc/tDhSDIrwnMbwAoB8LthbQ8FCX6MTgp
mDgDVfYOGA2JkRopQd6RgxAXRpD+FZh4GHrP0I5XZrs/P6WNU4TSoF4tBnlS1rVC
v9TW/CrYNkKdIE5e7hJc0zsiTSG3vPkHXzsl5Q9ZqhA0L/Mims1HgJLFGas/ijnZ
yxCtwzp7ITpYVhdsWSflZBV/gI9U+zXXcpRz2+35PVfmM9GZLlGrzAMm9iHgW5FM
vI41ykHqHD+Ms8lzVhsSGJsr2cxqIHiYAYml4FER7NNHEty8U174AsPTl2PdckTK
B8mnmMVq14GpO9xsY4TKVvMAJr47bBJjnfYHf/bBe0ItW9vRT5REMC1oMWghPH4b
7ervWuJetCuaVFOm5UdMDT8WHqlZq8yHkmgwpHXg68m8tnAIko0qfjPEptLe/acA
ZMN5HTAwtpiWpjEcKPyF0aqOthstDhmZBfhBrOzPaOzOqF7FcI/JLVxyrk7yNZnJ
BPudeMZfrDkvSE8pqd+CAXimN8rJyAU3b9N2+VODkSf+sWwCiX8xvZ8m7JU9WufP
W7HTUztXs9LUHyoDk7j1GpGJiacdRJADdUts5XkNj1TsdBiaSxMPdLXIPFEArNPM
40XRKvjXSyRLTRkCjY5BVC2g7GmWtA5LoNjBPBcQWUyCR/Uv/tUcwydhusew44q8
7W+YvNtkkN8+IptfbAbwdn6H8YDhD40KTUlPykdaAYJd00iF2Yu7qihzA7c0XldO
/+T8pSJBUvoqhFzTVPIDQ0SRUsoJfaDKV1Ct2IWUKmTyhoXWYRGR7sSYS7I9CA9e
7pxr+o5GEDitvhdcdvru1BXPp31PoxP5EMzy0wHP3in1Ftjnw40g9mcyn5ie/jmY
LPirLMWfzs/OWovAfREZnWA3NRxpN0Yb0kBbxPr96Sp55pD0Wqt2BQx6lYPAy7c9
XDKiKH/GGntrR2ZveNUJjIhORoQGdeyYpdKTWt6ACkWiI7P/HF6/QAYjEgkNLTvf
jkTgHQcwR1ZNdhxKLvUqghs1DDyKj/lA/em1lr/AFI6GdkrA4R3ymFsaWhyUOOy9
7m8aGxNtYz0vMOjWS8T/eEP7E9I97D0GKBtmuWTKWPXEjNJ0+rwanVkImc2iYujx
PuillIJQIe8Sna8vM9wkqUtn3JYkkuKxKN2rCBSU/u+3t8vaY4QboVz4cKsCZEYm
NFX05x5KYnMLtsTZc8n9dyOZ5GPcUW2Z3HPcodilZLBdJEJxoVFHzp0PTwjPi/ag
SxJVNAteju6z4D/Ogw9RC7il5+PM+h9oc2pZyYDiyROT5vaFEIUHdFc1EN7YufY0
NgbvvScszRnH09yUeaPnAUce7bxH4Fl4TgWS9fJl5tQBgVZReEimF+dMceXt1Rvc
v3n9MJOzZqIFba3da68DVa8kCEtqesejOCjfYezI3W8TwCWs5/OcnOYnC9VoXNMK
OTaSLFdK77DhM9r7ZSzSIHoWP26JrK32DKTZMJth8JatkkeXYjQK9Jy/2B5YZExx
XKPMtpbV/Wt2LPOZR0GtKzRiixRZKFF1NpKQYSTADKmEwbanP4i9OQy8Gr58mvps
Qv2R3frH/bEhoX7OumUP4TCjHdv6GCtEqJTPf6OrLZaeqySiEAkTWU/Owqoc5NlU
ezrTF7Xu9DRgYn8NJO9Ily6VglP6C2sAwLrelopFOOutwE9YzMnNNfqIXjR+OzkE
s6eIAtWz3MwUXSRCWMYl4TH4vpx8Z5WtpBEcSATP7+XI9Kmn2UOsfxm5QpJ+iP1A
F0XuXvmaI+BPYSpsKWv35yvZsDpwQbYLOPJpviYlUFnGUG5AP4XXBN37fqMoSlUZ
e7Gvq2e8+d6UJCIHnjmP77fQ03iC5rsOn8idvp4JymjHYd2z/qh94w+hQCoYMovo
hthkIOOjqwere2RmSQQ3OEIITJ0+DS77AmCnLRTKCbqTqvzinL4o9eJehZ4NUKYA
27yOASEyu0Lo28gjzswWJE7SMFCEtby7cthtAnXrgS0Tm4EzyKGCsDBp4ViolHU1
qQcKADAx1RdTmY7edk4rFOt+S5UI8ClR9cL+nvIK3Oor0QTYqxGVscHRDkU/GZ0X
TpZmyK244doHOR4BBn6y3tV9jAX1n5tz2ZBeVYP87UNoi1AM0QOALpQHhGAd08a3
ekhRRwvqtRzcPnFqlX+lCDE8RuLVgMFwD4pnmOWGIGwCvNboTyAKoXxMRuj9JS3i
b2t5ETlmwslZmCKKcy3tLUoNs+/dIKcvVaWx5y+tfJ8yXT6UtfoWxCey2p+0He7X
tjmG++4Cg9qXEiTMLKCM6LzGTWLkz0Lb4nBbDfARJoEPP9KOIctiJAgy1J07G2Eu
B2sQZnXDFNgxRRlo/emOlDxXQYlI8mUwMJdIfJRx99k8awp0S+GvkMPlErOQxbjF
5cNBhOM5vaIu4uOdzy9GXhIwT2Lfv6PVZRfxvFuLZuedHIFUxeJUq29kS4GlV2x4
D8FaPxGFlfyPGljIEt7dbYmlIwhMhqK/oK3Y3e7UWDPIFLkcXkcbILNQ4Pg5Devf
SGLxQXxS2JukUlD6ZObelhpiFSvH4rEXoy09minnVeFsjrZAN9IZ9PwFRkVh/Dgd
491MzzIf1HYCsn0l7M42Wtf7lsuGUzH9VhSfbP8qZXyUfBhpKvNVxi1o/z0TjX8e
4ocFRB6PMwOYSzJDS5RBTxxS+xyHvaD554EsIyfcnXuS9410T61W93GZzd4uOiXn
jc/7z6Jrsv3SGo4Ph/M6hP59+bKVw5PaQAWwOizfB5iLaXQDXppvvjUyygxBx1jF
CxI+QtS1ErUBBujIfBGrRGMXNmpld4En2eDJ67eYMisjeJlq02TX7fEtdQ1rMnxc
ps/tGse2+ONAPMq49pvkhuIuT9Kq2bcZXw0j1NYsi8QcDMuFeXeHmY+IejQygdZ6
RAYGHc2zbXZ5le+g9+eNMujDjksUeNPo2fPBaRc+kpoad42IUB7pTOqMOAwMKP5U
d4dmWAH/3oWGM8UhMfqP27e1ByNLn+7xMG0/IvjRnw59e+uGnM2L+6WkCztAhM9a
GRGO2OBB54vR4h1DZGe1gc8Eik/Elt+hWSqJny3d7R05atOfvdX/YuOWJ5kjpgiU
KmnAACg9oHhze62fiXIeHNORNgq1PM+br8vWElluL4hCWy6FOVWHGEWJrLjNOkDT
DtlL16yDl+wDLTYG0hrczynj+p30idVUrcUw6POs5ExjDmVnahoghbFElAB2e1I5
WNLl/J8ZRRlxgSa4/WXF03O5pKHh1blcB5vqMx2KYChQhxbDfNeYmC79TkYRznhv
JOZPW0z1pNUoIzMQQbMZr09lvlZHnQGqPeTciWbZBvBftT1yMCz6Iz44q+Kp8bjf
onWE/JKrBW9Q0cXqL5fXkAPnyd/zElQHLD5MfvBukHvPn1OSl91Uo0n2DnPVqdVN
VPJ11h0j/I0D1rLk0EXTqTTIksQuCzBvDJ/DiTcRciHdOpC0uNmGg2g5tPC03pyE
nFWVg6jbDz0wCFeFVyGc6eatJOTW7VSEvob9u4dQt8lYbI1/Ejfs47N/fhHVYfP6
BCQCeYCZeFj5n+bGDWR2n8tm20bYzv3gSY4jTG7izg9N5DGeMbSfDBBQBm5PnqbK
RylTD5b+mILla4qC2xSL75G4B67N95zL8nnqZLcK02agxWrGSsYggeyALXa3ZZA4
QwzkCy6JQb8pGYBGcNNSPAPTZNYCqrQ+0SzrE3cfWmpalfjFXg8M5Dm9ueFPR/8I
os0KfQLFbkzHyoZ7Q+CBZCvftEU8DKjGOndLNW+tg6PKmAdtqEE12Io8Fi7s7s/V
3pWbp10deDB9SrfZ2es3MttooMExErWecO7TdVhdAuGCWYeW7d3Td0xV5MOc3fzc
BTFGPlYtT4htcNuaHlCzgYicUc7ff8Dync+OBaOjbwaLLSdtArrsAgC0Kfg3m9X0
E+5gJn4q8XIG5V9tGmpgeY/YDLoYCB2kdy04MVqVKTPKon0rk0+XD4EXBbH4MPDz
vBAIVN7GVL1ayP3m7i2PLAohvRnbErKePqxbU/DeG1uIJVAaHBqkcL7jgUhKtJ4h
w4fW9RShKQI+7Ra+xfL3JiVXwKEN4ODZk7J/GhHg9+jLpqV1x8wMwvLf211wCTf4
bGWhcJgvnvvms8r255Jng4YCqAWgW2mnG59OifXopPECAnWVRT9/rD8LsVzYqnTY
qwWCn0T9ix8ZbtrxghPtOM1yJmkFEZjkLP05cFaWskw0XV65mC/O1IjwscIsqb9X
Cqzqsb8bXvJDzjdlTEqBLykNqisvUpKoGYLVivqOfRDaXjfTzmkdruFSKg/Kp31R
4MrPt3EZoE0r0X1PlRUyCgiDyZrtyS2ZVOGdFIrS13yeIFl5fAO1NzwaKUOBKN61
HwsMAH9dH5Q6kH1RPA3WaLg3IBYfYyvLd0wPtEyFIEqpnGuMzDRNylspiyEAGymP
CQvPdG8T4iT1beLk6DWWqtQ3fyRcjsaQqtVkcQDzLf2nhK3DbctM+36CCn/mk1iR
ZEcRNawMsU1UpfY3zwljtB6J39WbSLwJktUzDMWCDMhTZY3IMSKoavHvOh2r87mS
GqPgWabl92iaoXmrJfsOD8f17H3KDx3cPoBugHjz2jxfcIpKS+CW1f8R44lhLe/u
EAwtOM84ZJQoRaSG8LNBInWPsB/dd583T7jmWzyXOfbwPQ7npgo8BtmY4NZIsmS/
Q63Mt1awPdU8fGCXo0uYFGHu2OP33iTmni9tyH3V8ix2y0PH9yhLcMxyYbO/sBAK
vAhWGaAPVXE/nXLQTUCJ1FWbPOuF+yICe7mPpsWnu7ud+HlnnZ/oDFQgjdbYyW1J
4O9lKDUrBqfL0yjZ2ro+fiOuvq3DhyHFWiKm/0U4b3L13jj/PrG0anasl+sUxB3D
5+QrvIV71+O7jrEgS5ti8aZlvNRocRwJ4vKr67VYGeqwM52SoML/CQHGUUVn8Nsw
DKKFQhGD4+D6pNnkbORcWsHGf7oLdlAQGW4/fPtGG07CrcDGDz0pW6kEEOSQRQfu
ceouD3IlVUDyLuf6u6TEtHCHEdulLCRf296gRhB7u9OKZkh6e9K0tom6bkJpiyS9
nrgRzClk923GQfERGutj7GdnMZmhzv/0QNs+F9d6yXo9ImIqwBT504kASnGwCPXx
DkTO7duhkyeesvKoCFuIANVhuJBmvJ+02LA5Ur0QMZy+uM5T15TeQidb23uaQlDc
P04tVZP0+utkOJ78+m60CtvYHmU+9JTSXtya7QRRHVN4aS5hF0m1v/XK0lrStHt5
+nsXG8TtSjrQub4vW+BMueHj2rm6OPusf9mJgDvDPAI1iJujdiB2AcEKh73MojnW
SVmJw+q5irKa/STw/vud826a0MCSv0LLcqZeeNzU7X734uFInxg+NbH1a5eXBXh9
5gPFxW9wAR8shyT3AaNjTxR7fRtTpi3qwPFOC+Rr1geSnkv8Y5bJxGw+jgpYClqP
g6lFK02tuELY7q3KCfKVZ8ZC0TwrL46VSTab5diZNvA1L0mnzxjh/eY+VN1dAdmH
t8dVKvS6BY7SHpGBi0waEHIxwR0kAF5Th1l5ANWYhwdtBS75hHqX2kGcren2/1yY
7qiSa2kw8cJ0qwPv8BaOkdSqYlQcII2cLq1a+BOIgTklEHolYgJVHgo+cYUXOR0R
fEqzbrVH3oAyC3SrG/So6OgTS0dj8O6+o76dy1jlGR7MQcl+j2nIa2J/s+z4fbnZ
EwuFZpEoQoc2YGYUDCer4peNnlGb0wYpbMQyXxitIRbniZkrkURUXT/3AhK4aD99
ZMFhgcldDZToEH5jzjlWxfMM+E6HOz+od4oxdDCmVfyiLfjKa7cc6304bUinyVEe
Cr4qEkSR09fmd+VgcPYlUBv7ogvyirofOLMkA2EJDvap1I43u+3yXumrudC8aQHR
ZlRF5TK+VjcnsKaBisJbZgJZ9TB7PHg+4NO7ZgsTpL/OOBwufdengvGTeOWHKKRE
f2r0rVDaaQUwxCyr0gs1dVwnB7wd+LRS8nXL60F+2T7kJJwqasZVcHXxn/5R3Y+3
WccBI1GTL2HQFNn85RVexvS7ZuSgfEeUUHQDvh15GxFruR3SJvH9qGUNGX1yMJP+
EmdyEmh/C4hmVF6F+kTpM+a2WIu8TJ1SEFevZ5/9E8Qh00QkmHiRx/wRJeY7VdMM
pDnuU5jqqzoWjgfmbw6C+27xzUNicvn+ACqytR3CHb7Ts/G8EJ7fQsNnhszolLGE
CKYR98KCuJyjgbulO43wMUU4mCQiQ/j9hBNeIhQyjcmZF06cXPaJnLrI3qNJYAwy
t4CyY+DTqWYgVoOdw59XDcSLmGzMiAEXMoQsabQEC7RzOVm5bROAOu18bDEiB/O5
Fqr76yM54q3WV8buj6DhhScCSHidRi8qbQDqaUmmH3xPGbLZvUJbTjx86dZ+cD8t
7AYy2nisO+DCt+JQNgFPrxKqyIgjdYJ3ZZTdwBVhMqx7fhVpW88pVxb23rr2tQPF
A22uc3ux9AQpnBe0qAET8JFADbJlcnh2KUs29pq+r2PKRwXkh0/JnD1Kih8kFoyG
kxkTWS/eLZuytvtcyB1mNZJxGiFo+hQKdY93Ug6V6HHi92SW0Wl/x/WRuAGlg4fj
Io10bW9ZG91tNRQjquLENmbI1UwbKAYlwrLVBmMFFuY4psQi/JgvC6pJl3E+q66c
Nh7InAQ1PlTW/rAL5QZS8kjNkUHmB7dbodkW0TbsCzYnz57Z+klXPLOkALYmdwRv
laG53al+byTnBFZaags3U3eNER4cUr2HhHaq6wkJjRN2Zmfj/zuRuH7VHFicoIXV
okOAcuKWQyUJpMw0pYWN1BLmLTnFwKl+FjhY0lEA0NAIA6mGj/ZunwcFyts6V8G9
H/caNGbV73tKSAgrkz1pS+wO+GKSOenAypa8aENrMPmeLMcnX9fFAXa2ElYDOUKU
LtWlKQWr+hy0/D2H/0yZfDbybLv7ZoMXhj8uRsZyozU=
`pragma protect end_protected
