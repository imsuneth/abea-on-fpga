// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:54 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gA3SZnoSvtqp2Q7ZKz6pqqtQLaSpsxlCOVfaZglD0MGBxKmQbkZZvN/3X4yuoRDc
xm3NWfzlJm6uKKEo2qVSnJcaNFpVVX/WMTrQMM8xojcmzY6zWrkwgGHJRiH4Z62O
EJAwLoEFRhUucviJUVYQ1kWzIt4ysoStMh1qQGUnlF4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7152)
sXPY5Fe7MOUYoZajRQcUaxH5KClepP+qLd/+GPOfn/lbpkgQHuhgFlkKnHsaY2Xs
Y6ehjVuDD4Pgq2s21tUdEYDXAvt3Gi0lR/M90g+KQ5PiGbIaGoT9FpnndgNS71Vh
la53dM0Kgw7gp0yenhyfP+xPgB5Zjfr5ziTYzOfP/al+sQZ998Nt8v7kEVaQ32KA
Q4Eg1hQSmapa2iVlDrg03vp2BCZMT8xObgb/8JZjYyX2cRarXZ/LXXtR4i9C2W+Y
9pRwObCdJawD+IHa1AVc3ZlGGCxippRdRrD8tA1Pey91pWwCQXW+3Pwt3lSQ2r3h
s23bQ/lKy3km+4iY4g+QkS806hIE4jmTmF2V/k2HVS/t0kW+DGLuJIbLxwIG0Y73
TNns5BZbz3HWENgNtFvhw/EXvhJkbRBusB3yRwpkBnnQ9AhBzhmWQVFw1RRl9wcW
/5NQ14cjsVKblV+wahPY6PL+UoSOsxKGGP3I+c5MQHUJCsaBvgNxHAFZon7gbYks
xTz/RM0TyX9y++y1TV/brU9uxSIKpgXyUzfzPexR6u24XQaijkZsVdqri6TLx31Y
fCFxHi3Cdnl0X0hzIwa+cRzQoDNJ1SIksoyYM9jT0HwQQ5+UBdIL9YoFO5qYuhF9
YUoQO6hola2IeUD2f9rxC7mxjCdjvkfyqJoMdpt0r7YCfM55xICf6h1nhcqsg0mo
Apa+aoKyGpmTmNFrQrxu7YxqpbSq6xSinl5vrHr2AIbijgB1chr11y4dNKZDeI2M
kB17sr/5zBDDQY3UHUvBnVI7+w4uaRAS7dq/EG8cBM3CCmSbJJCqcovWBGEI5hSL
ilv7MLM5zH1F5X7oBemess7Ashkxc8aBPvrYytJ5ax0BKZQNCFKIW0asxMqQSwti
qyJRbdl/h3oDz94rnLW0jumdKLr9yWCPR/x8XMl1MyFy91964tSrgotRtJvbdLFZ
K80OE9jUuQx43E16pty5CYOj06eBp152DnB5E6bgt0dFDNJTVPYq6Ru1Jy0UC0Tt
35wMR/wxQZS2aqxTiCrVhXcbplE2uI5X5BWsEAyI+e+4BWlGilwyrUzpafNSsSAt
AdvyroMBC9A6j/LmYb2iUFz9I2sAZJk32bLh9h848iQklIFapMN41IXCepPJdWwP
P+sAPQqnv6F5uF58tjRHV2KdToXteQ78L1ow22c29gEV24ZCNcC/5SFRdEVC7eC0
zkONZN/S2qRrfmXKRZkep2JQ+t+CMXZPPfKcAh7JaoSObx5KkCwxMb+Mj6lrmu/z
vtJK82ZEcXeO3pXy02te5mEnLzuN/qKa5GC+HoGvL1+TMmmblbm1QldQmXWnKYgE
M6m/UCOslAJ8Uk7pRBYwEjuLY4oF/jP2gs7mhdMrKoAb74WNsqrgcxtl54HTN/gO
eVy/YY9KTlyNFBotkmEtGLIioq9eOMTJB+PS+1rcCbw7g/cbaqOGG0EbscX+G1fL
bSMYYAJxviRUotNJmbU/6CcUo+J9zIyKofBr6jDjQJfroqbWbtMRKEsvR6DQvq5c
AQAbK/FdH6XB3rIb1eVUaloaZxB0vYk2voBL0y87hNKjt3PhWjA7rNCzpncHS46f
EqBBIjt+FQyeK6FdpT1zZvOLIvb8IgM1Ge3SphgXVtqoZSAEY5yoXtpoANi3uY8R
9pDlbCihByUNPN7K77gwUjRnb+A/ZYf6e5JK/7MqSHY5UVKOOnQVER3D6cnUO+lR
eu5jPhHz7Ptexzpx6GVe9h21I58x3W+Xt+rZaNN8vx7uMJuO/BzybzZXsrpCozu5
8htXWhZqtanlnwZsdLd0F7HrLFy3uMWSgxQwBbxpDbLIkiliNeS+CcstqOlsybIA
XIhijBEE6OzV5uRrHQtHk3u2BoqUH6PdJDaXytF0sc7WdukBIMc7y6Ss0WQP1Du4
BW/JOsSyaj9CPutsGZIMOMsrzIa69NBcgJVcTwj/vnT9XTB8fGjLdmFwR2wq6JxT
WhclA26gMImcNm7evM5DLUh8C3g7L3r3oe7nB7wcfvvD5lYnTnf420dacnWmqNH0
yTpbB9VlSawwvrd76/powoAUEG9S5r2BeEOoMtNRFhmzQq840VkZgqEXNsK018dc
bQUqw2FD5K7HN+zbm7Y3LSwhJ95p2WK09DImC1l5fxrZdZ0+CuLEelO4A0PYHX/v
+k5VutEjzQkRHqrIqgrv7z1Mr+BejEr3s/mM1gSHh4+QAiy9Dc4SN6EiVp2TCCBc
XVzgJ0LYO5iBfUjy7L7KV/vkh3uGL2EReK3oeczc/B4C8sCpNOnC59MV4r9q90WK
jiYVSNgHafFi8Z5xCwQVuJqHdqNJBiPiH4z0GgMAubu69RFkzTVm3GuPbCW2ATp/
b1TKeAnfeiJuqT5WMRdx2P2X9+pqI4iSKihJYcjI2VVi+w//KCr7VFeqmg8OBKNA
RpkV5WJ9LvvYC0OdwYAHqMcXW0of8m3KkKssHf+JRz8ZoEUL9oEOhKauMzMdyGHd
SEOzUB5M9UMyN5Zd4y2ooJiZzwdwGNMZ7DAOE65Xaa4LvZPPNQqJmyWUWNBax94c
qp5ervTw/2tuevEESSx512wiDXQywdRooIJuYLXLNaku48DARS+5DFE/FOgeod/A
2MdLBU3nwSajTGpjyBFMwZZyHxjQHW5Uu1yGUN++El8yvGyFLfDA1nOKWJRSYgsK
QqIFfePx5K66PoCjUBYlJxeksfTW4oHFTPt5qOsKFvPJyDo29uKgWBxEy+jOB1gc
2Ro3mM1MSSnt4ShxCPtpczGOVGRHqhoVdqZeudmEEdABAwdi5NiA0+EY0gI17DVm
ZxWo5MF00DhbDVOdWUWJ0Gy845Nv81be79+uxlwy4tg7XMIciHOl1wBUzPA80bQT
9q67XC3+1ZTXXJXDhF+QzlyKmePpgwyUrrrG4FcO494QzgMLnZ8zo4V2xVkiHL+r
QTKZWXAxkTNihUwIPvG6WkpMGFM46v0sErL0Vd+I0xV9rT5qyHSjxJK+ueKIGsls
dOEvIYv5uWvywWNsQGNUR4fZwfK17EMOfoMUXCBgU26YigZxKYG/Op6r+gF9PJGk
q0F/APvl0lLSc2NJ6350sAOJAbOTpMLH7jglQav8SngpPVy9hflkvGNcXrGSDZCe
Z6QE1M/xM4ne2bjlZ1j3c/uAm63QIBL6snX5tp7X+hHCgsYLEI4VL7s/ayJzUt5X
vr0/iyAfpwC0V/9dUDq1H03ESDbaS+XGW6gQWWvOY8RF3pqy8aksP6OZV/kPsun9
0PyEpjeoa6q3Rga5GX1Y7IivQGlhJu6EHX3IDURrbAiqCvaOnYHWyqAuX01LZ3t7
N8DD1VjcO+oKriGzNNYSqso3YUWJDr+MqRMt9GmIQOR8HoI2VSmSEWhXYdsWsIJ6
8u5+qhE7U+LUairv593oIrjUsNwe2fc/jPTtCJPE3PT+Tanj2/bWRr3C+RcdZt4v
w/FETaXV4AnNrEGiWXQQ4eDk97KFaG78wK4kve1LbjDWeBOIfULolBVrB336AiDn
188iNwZ6kN3osTsTPYQLWKa20miUrc4KZ9ni1Jt2e05+4XKTJjP0rQwF1Vd+FSxh
F6QPEroI7eES/USeqsh9BaZ8+tsjXfv1JSHbE1LJc/qEYeMORmus3sSykLfJJgNu
dVKTKG3ELrOHT2kGpKnirPblcYlNGU1rAWjCNti8hJYtmfMNk+swKwqlKO9bLGQZ
fkncKmkWrk8GOaDVzLRTQ8IjoHulX54HynbkGtLbBZo7TMPl4IwNsMQTCzt54Icn
ML8+mbjf7DEcqCMdo4xlXbQ9IMb2PUuxuc8gR1B1FHHOvqL6p/msAFv58MP13LtJ
qDOUk0UTuVHMkZwcKCL3dgb7gKHZt2yEpL/h1B0OMWe9ly1WP3cpr5ErZTgD37yn
voozw8slWgamaXgDd8dH5GSf4j6Ln0W+W/bkQupO/uZ4yo9bdWcCXt4Qp+dhUWrz
PLYBkbRDuTyT+Vcnent5BzX5+/tJ9sikWubBYTKFIvUVMy/0fLcVdVREuHeZFomy
DVJM9ohawTR60BE90/Ev9SwRytXO9+mb/HtUNf8de/6De3zA0gMQVae81LiYD8Ds
UallKfWGFrStBtvfeq2tlTKRoAOUhf/cKwdwgY0UDQRTMcrzxLN5bbVta0OUbxBn
GyBHiNSwjCjC+lhVZz40l5jiJINsh9V1Xm7LL8aBOQ9vEnk6aBqDsiUIIWTfRPGU
0s0h25xAFeOGp2lrWB5jnWuzmlSDLtM50mVsuUadrrCydSYoLqpiTcFASmaLizye
xmN8X0q83jddmt9rFW3ZKkWszLOdPQCd25S1CCCvVsMg1zK3jMHC1+MF42FKBwS8
r7JbazaRIxnFTZAimbSATYzGuuGhNYrr9lkhef2vNK2JCaWoOugNomFP53AHUh2J
6E7PjKXsrwsp0aeQSim09zEkCJAQeuQCW5MBvW4d4cgn63/Z3gKSHAfX9CIKBNcq
HQOuCFBU2nNTN/BZX/sKcAbAx7/Y1uqvg/OZLQCOErGJ9LK902M//fW4hxqSPRXn
X7UKw21P9r5+bMjXtwYfhicdhUelzataTqTuH/XDxy9K3OKjPa6Z5GzzKQbx1YcC
ogDWnjAFkTDD5Rm8XqzezLki45/sLNTEkhpZRX/yZ58ElukKVh9FHFJfZrQrptnS
1BmZ+aXlaGFJ7LFcMTFX2CQkwCspZJLRi01u1O5vLYlzsLbyhLwDa2emDlt6eyKc
Fr+uYV1UPNO0Ij4FcHtMnmY15bgsiT6cAIa8EulDpVgIXzQVYJ7O+q60kyLpeIEA
q3XU+1A7/yURpq4lpWZMvcq+NGPgUGQm7eA/vQSuCYrRuspm6okuZWaPNN4mIYKF
z6E19yLNCDn5wpzZgnmArrL7hV2KHyWZNdGrWSvmSJOtTH6IMVyHjvysSVd30wFb
n9iB0d7jovOnrvauCvm6lFyKR7nuA77+c342QY13W3Ud+UawwkLm7wQhRXn8aFFp
S4REz8QmN7zVuSoFE0V7OFQrtrIVOzgDLNpX4pKrrGZNh82bC+knSCEV50k8qpSB
Ty7gGsyyG4LcyilEH/Q9uTfXScncbAtKbuSml5BAz6tVeeAN5ezdpYa+c9nyzILS
x7luajKYSGdy4XlD9cVgN+wlUP6vC8bZIHdM/9Dg8qwW6sglXDGCCZ4PsRLJYt4o
Ykj/MkS17a6YPMXVqWDw+yCQfnRZdns5h1/NejuYYCFEANFq448Ox8DsaO4Yg6RX
NTYVZwlc/M65Cb/VSbQVo5r1ZLDLGAf7CNSXXand/EWj9Xb/NZC6/EUjXZ3k0FgQ
xx5p25lFe9DG+7+5uwijKx60S6IyxSKb3i1HQxux87qPKqgz48wekOp6SaQwY9oc
xdqkp+hQP3ItlReVXwrb6RwqhwPbSyn+HcrFVBS0D1wjOLoWgYrvz2Neif09vueO
VHHHCDOMHfqnd0F1yWqZn8GnNRx63gRGZv/S7LOFuzq7Kd+F1iBHbURYjb/hYGjp
jllAuXjz7bli8LiPTezJoXRVsSJLS1NfgR6qvS4OSSpYf/H2kHkCzgNOIQ2zbpE4
rNnXz8ov/7b8M/C2PgugSyK/Twa9XfCHLP0MWzy2z0KKTef7hxZB1ljlTYRfe4TT
eEb0qpD68oPxFLKon8Fg+CMkOku43zl0zLOB7CvATytFlhz4ROdFcUOTCUY+KtE7
hP9a86dtjBZsDvYLFzgaEyhDEqYpO+vDwz6gFoo5BNKcZqDQwrdyyigjPFR+JzaS
KijGWgWZeaiKXhvPwH8K1P+1vahF3RoNMGSO+vzOINUDDWjmeM1keQz+NEUY8I06
dSaZvVmGh3lsrJtp+cIxgmq8uGzhxMVNB/PtUzFfaYtT5zQdmjMDaWYtNaLvGA4i
cnqagRur3fR3ANoi51xRjvV5CZ1QBRuSBNHpM0/Oksk4lBrPOiz9eOK1SUMcPsHE
+bw1v8bxAbO0QlsI1N+muRtqStvbFKRh47z8CU/C4oITOCS3b2ufyrU6DGXiwtF5
iK5vYcmuL2w+WcHvqHLKL2kpAqCCAJhrdOoYeglRtL5/ardbxOkpliNRh58Memfo
uPyQbwg/UtFfwuk2TqB1G6Zye9hKW/l50YwEGN4DZDL2aD2WxIhWyVrMOnQ+jA60
5Bzurwc/o74BToO1v9EpEOymEB+xTOtCE7clppnA5M88EzrzLUF2nEEUzBopNyal
v0FbK3/V0WmcSmLGAu1QNpyS9ZFh8aV6yrvXk7d4jKjQXnbaeTJrJSvN2qesoZ8e
gh2eJco0sDstWVy4lGHzdiw1y/oErJdEQrm6QuRWsFAMdGpUpo+BZ5Pg14B/zbJZ
mUgkPWRYhrv+PjAmgp4v5/GIlFEs3vE+JTeSdrx1P2Enj8pxqn3rD51gGLSJO3pb
AgCVN6FU4DLkDFFoA1NB8QhdcuzEvqvFU6dudLavbpyYxqOFMxVS+E1untIPl9C6
vS2h/exMtsEGCdEiHfhDCbDp5LME1rOikNxdHJjHim2ymOVq67XE+Ag3rkP992JO
OgQh6D2EjUHgh+yv69X6zwOiFQIkAMom6V1eF6gmFD9YVWXy1QqzwhT9V7Cm+s2n
ydTdrp5u0h0/icAcXDw+uFboQqUCCQXYM3Vp1TuEx2+5+QmAzzpzNjGhfpqGz5zX
WSeDG9StWAqVYmMCXlGsXrjJwx3b2GsbTrmyV0toQteiRDcdwknU7ymn03NI7f0v
mNCxPSsIjSqswcwRm4lAvyWkgXUflZG4lE27mcukoFECtAFFPgSTdVUvFgSJTJXy
qQ2bnA1KS+FvhGRhzCD1ce+w8Dm5iW8C2kGGsukJTroBo1R/IhnIum5e2oZ9U4Oa
pJiJN8i4OsYjgBMTGNaPvZdPIcNj4EMmcBtRtehEYFvHwfscQHxeikORY7O8cbIQ
mBIZXZQokWeVydSgNbP71MRNeTBll2Q6K56saTpEjF7TrY0TXX7z6B2GPR05/kH1
mILZ6I31jXfr58xr12hZS+bWXH5+uarmQumO8ksD3oZXSX6m5N/m3Ay4x97Me6Sn
nXArV0i+CN74IaTyqUcxlKVJQCKxG28UJmHoAWAObtH9FQ4k2Kmir1Ip1TCefHZi
2ZTK48vFts/TC+++HsRHyLAM6HLPcdR0G4szafz51Xh9TUoXfxHf178fRElScBbv
wiebD1MwDzA/Hj8HKWTedFjv7JXm0wDCk63mjqXPEWpCMlTSigqTJfPsyKifAemF
uQORn/9WE1HWey+Ev0OxUnLzRMFa/FDkqHNgSxk0Z/aSHgPbXo4Q8eSORsvZ+rfb
j4ooRjWFU9I8jKgvFkL4LhiMOcyFeBgHTU5KrbYqaadm3LDwsLwgdGJkTYIEDCDL
0lXp60SZlnf2YO5nr1SyAROvj6pxwco1CuzDIsimQfMdAaKqbt9Aq5Xj18BJy9ZM
71p6fsocg121HJJEr+FXmKyHq+RUBZQbKdhwNHx+/ake/WYlKZ298yLzecFjQZMa
oE/KKGEiE7XEVytEepkPDoED8GdCVblFABRiVQorS7cJfvG6wEeFFu3ZsyaE1G8E
4/9mdHfMIL/ZOMRmkJevt4ib3EUvfxok8cuhoncqBqP7AwEM09JUgshXd4dwOYlm
7cEpLQmK85CmC8eieOShYSj7EPDvFYQxJemOtPCX6CI5PhxDzCEsOwieFBOKRvOa
t5ro2SZe4qyS5lgp/JU9JwdGI3eMCIQa90jvg11n6wWok+4ZDBbPTJEGGwqwAaqZ
hb0cT+ThwLpwGyQBALn6xg2HuHskkL9yHFeEO8b9t0VITipMLAKYNo+Tyaoi52qY
TLUQhzc4Bg7tr6QpLLFUdZhIjQD9LmP8UWv9ae5lYeefBx4L4XTMbxpkWL3EHCc3
ptHG4Ao+5Y4lUu4VVWuQSMwYMB+k2WfKwHZeLhy2hh8x0SNy7B4Pkn/xvJqR+P3B
TtV0ZWAri/y3RL8nmkSw/hprW8rq9WM4DGpjLWhJrXpsdDkZa6qqCeyAvjoXBhLY
Faq2yZL/JfRS6tzWZIn/FYei+h43fNUNGETQAdctTrKSrLeqC9BN7NfsR3Z5MIGO
HtSu9fBf11pkzDleBpJP7Epr16B7VnKxEYoj+fkKaW9LDHTCXSbBNiSq6MSh0gob
vkZLE+xSdgSCKlQORRg0/jMOfb4Zj1GAPVimlw2VCDDPoJ043f0NrHYxOV3foxFx
sCe0GaZ+6MRRuEWhdVcIEmoTbYuhtXLG/LdmUGfbV2wObX9V5uCdBjETdJR6H7qt
sA0hnmv5KFFOzCqRaMcQp6DwkTIbABzsfCMMg90Hwcbz2cMqdPXr7Bbl+DfsnXq6
Il7AXubKIrN9WUi7gzfCgqLItbN5m0F6Vk6JQQZJybxQXc+nGjVhaSG70xtnX6DI
vjdL/J+YXmLjcRcfekV5zT57kJjrB2wSaTleXIEfCxzkk5kvmQqsB0J4NoXwa6yW
LjvMKFIuXzPDP9R7OUs3gEgFLlahVEz0chEMGEGwX7YUzK0UtImdcmzs6MitEnYX
kFX1D0wL6MrVogYLCDHwaVATebkwVaIOLP2O4hHVtGIdzNZbWTT9Fuu1rH2CVcwo
tAMnO9EfyZIIOKnnIKKu8hg7EzXT6nqEiK93lBDMUS1anxe5/nz+g+WqU0NrC+60
EdjFHBqnPFeX7kZm4eC1MiBJTIgceXRDAkVZJWa7lNPJ8GbG0Lqe65Pb9xyULzxT
b06yMytNysYRN7xdXWTe4ttb+5nRk2sWwgCodxn2wKw9sp0Fv3oituDQdk9rX108
3AOnjeel2Anx89CKu5RVFHlC+2XLb4mqJ896Gt+zO7JReFF3+Fuv+zkld3kXoq9E
9TJt16NRtfvoyoxAhHROjkJx7WZceLgBwFo0CI2/jAv+RRSsnkqyM99uxDhhSxqq
w2gsvn3N4bvHIjNHmFUu545qkRFGPsgT6nWLLk+72xXLVL/DfV+9Majj5IlZjoph
l4N8ut6vl43HliZL3imEu1Kt8ZkuatxIe+J8m5eqZjCU/ugzdbA1J1LcELRugqVw
amt+OB4FxWkJdc9MX7REReH750w6ZNyaVqiiM8jIMEL37jRVUosrOWStQhAoIJ2L
xKxLQNi0ET/JzKtdNUuBi/npNR2woxiREfXa5FVm/11tKbm1ZZbOqssJp9JgT0Mx
aPpTCVTV1PamPVyVpvplqjRQKVzc4EOv17CHlU0P7G+Ow9NKiMLZw0XaTOaYHLZK
SAHopy9bdgRhJn0W0cUWexM1hgLTzL6rmLZpNjwbjTuuG2qLd+X83OJW/3v4PUbi
x8QiUwnsvt9WbS/reGO3gmvteFvkGfM2vmz3i5BZMYnq2RKECXfBIRN8jCRfMQsf
4lgRl7X4pELiLlLgOMEvyPdCNZdDypLLGmILXguspQS8gQv5D0CIztcIB2cQ3B8+
g0bHne+i+puPFWhMSxV8ZPUxrtRtWqyRT4AkpScNMlenIGrb/lM2SDqyA330lMR+
gm9VoBlrbSnt63Sk1y4JbCGRtRV/BnxMwav2+1fIkdCDBCKbgiBAnILP9eH9uTxZ
`pragma protect end_protected
