// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:30 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j2WUacxGX7Z3CzYheKFuoG0LXlhEt+CRWofZfAtvTNPF7Ba704ogzGEsLtGtSmdV
SlSmyl5wfZuDp3I6KkgDEmppfdnyIeD/AwYX8BjMaPio7H5jhvp95qnS++CbyGGu
0aVJRalBpleu7J7Zym9qDBCGkwUk1FY7NGVk7NXnFoU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5648)
HSYZGqC+4ATiOo50g452Y1lUMnYV+o6iKCqKCBa1UTneS2lY/cZFsGXJV/IhKDyQ
jcE1ASXX1nUv6N4kBbTB+wkhdDAQz683ue7yVKsQ6SxiNpePTKh3svdV8Oepy+HI
vXrxXjrwqvVnKZlH6kAt9fiULYLXt+XfXjna3Lz6qQvl5+pxY3YjIC7bHY1D7MFf
aHkl6fPxuTHJVKz0bN+bgyF8sEuBwZyUgfNE1qQZ286I94Kt9nYp8/LExbPJM7G2
kYjSapVrqCC1C+XrkROuz9GiL+2xBIhiU+eyW/IgjpTc3fz4+eCE8C8/f32EuvZD
ppHkLt/Z85cu77bu1+wRN8z6aegD0lbYsdx+JztwEd2x5IXO9ZfhIA7nzZhf2QOG
Tted4Q/m+4lYePiG+abSlWwgeG9QDxVZWfvrFnoPQkoEq+j3jaC7B+Ch5vxFFpCT
QsbAltG5P/WrtEXbqri2W82NL1eHZQs03oAsVIwDB0TDCTE+ahb6A7QPLBGBHU7N
bTDGNDMfTRIJX52nQIcpUUCTjRmyFqzLv6a/IjHtvk3RR16tIVKrA2rMomK6VpJt
GBDR9kCJgD69cO7JIHHL88V5N4u/rwglvFxkqMpJtPDQ2/jynCHEKcAMoNJt7TBd
MlWuXZ4FJs2rLpRPeO8HJvfp1kSrNA+LyJnJ1QbtNZTT/gMp0uUJAn8zbY1Llx9c
YQKojmyoEHlWiGioe6kg2tKxyOv3vVWf6RwIA1QfqYcaL572RXJyqYOpaA2D3+I4
ozjhE44VkSHLs4YR8VIkCbqGAfC9/BTcO7/toUDb/EGnNeZL+zfaDIPuZhwmNG7v
Ysp1Md44+Hp9u4OZ4jDHkFgDpfqDv/+fzjAmgf3itmCmuKhW0VmGVksse2iKWaki
GjxBSBncvliOBIlbkwhlYQfwm0ABXYb27X815ayumwv9gEJdBk2y4+I8E8Q8Kxlj
3jKq1BskH5/ob1mgg0HngtY82XY8UKphSwxlBRAWZTZwWpe1GXcjJUjxSjAKfeDY
nzvuJJGluOGtDMQ9t3hMVYFJfGirVWG3AOTt2dyfW2K+mVs1pDWzkSs0oYZp9JZI
udnuCU/x/f/5jvm6IEH9b1j9dodXuOSrEug1ZFLTGqYieMGyrpQflKesf+fXMmjw
ZRV/AQbEPvxbm2YNY8636Dt+THaFOd72GrJT7i07vtB2va8MN2Efai5muBg9C38S
d0Y6yRsu1Wt3Yfr8ACt+naQXT2AJ1WI4BDYJDKjyVIoDVoOXfat/hKObDCJLDmUO
CdnydjqovlQWE7ymqa2ZgauAlpoBlNPTFAntejF2TuNQtkfB2JKINVzFyEBu5edT
tFAPFGtJanKyKW7oL3aeHPRE6o1GxxhJD1gil8lX+vrJ0bWiXMwxkmR5HbwT7BsS
eymLw4nrfmFlR+aKt9Us/C90O5NExSgeddp5yZ9D3Ny4EWfpmfamXVo1M66l9R5V
ApgnRfU2RzlB7jcCNz4WDn7wFaQX478fWxtOtATpqXcU6vcOYkXWWhAmbr/LUOMM
GAs+S9VB+0+N8oK5TPoPttxaAu6/6rzHscA3lax1b3YOdv7K8Dt7GfET19LnDhKS
2wWcSCbfnORQd3wbIAEGGLnYs4rSO2GBzRljfcVbqig7rUFnnP4elsBDrCW9IUHY
k+e5Hp+2ZN2+8YVJECcYKqEAk9T4kq4AcBfKk8IKK4o+azT5ENExvy0BQQdq0o7h
8DgKjQW2bDSPPrfo/DbIGTG+p1LENlTVi7lRyXTqlY7H4m80CFwCfk59+gZUfDs3
3bURictc3+5mmVOtDY4tfvqGfkqyGchpBtL00ThJVzF0Vk8Y4MqC3ImgGhw0wOv0
HqVrVjqEB/UTqRw8Zdnimb2i8dhbdKyW7Zc5c5EmRmkGNRQ+HQVKETZLNOhTXmTL
4vLVNye5inevJlSud10g4ha9U3Woke+rj7dQrEiUThzqMFOoe9+8XRIobYqf1epo
WJ0U6b4xYHWyni2LLKw8u75x/JfhbPXqrGH8F85iYrXmN6RvNPaFzD0NJ8L39cSq
Q2jVTXo6rlkSA0qpLBaT70kJsTJHp/RPMkdYntS5OnV6OeJejPdh/9w4C2SpwdmY
WoJONSbCZ8dkAd8iI8b11GdKNJlyz/0yW7NfQ6IxXEJuklbDoyxBveDdSAcmQNIz
M4dEKcSIw03YMuZl5cQhgQ3malLxkAdmqmVcZV+EWf9+73MKF8qL5CNZDxfj0IT6
L16/uqT7h/dWa+e2Ffl+ZbE+ZfdrDKhIqhHBusolKj4AFSslZrRoi81uHLZ6Enap
BIfSGBhboFYyTxJA+m+ocpatth5tJlpZWZzqqfYuab8pWxSvldxDZDv7PQEaYpMY
cn0WAjAYawwjQDvSv8Aum8w4X/bBsokGUjLR3eQWk/kP6uZlEXH02+qgCuDNp4MN
3RNPn28Xp00AD0M6zJnod1RqTUTaqMoYcKx0VIETQo/SDDw6R02+YYdTXdROpT6Q
R4Bwgh/YNKkU/s9vpwI5W2GDGsazCuGd84G7I/BXQKRIRYvwb837BVqHZBqnmvPG
l8H7xGtG6kRg1Z19fPUR6rEPOwnAsVOaGBSAmMdIvZivelnVSW3JNJAcJbm36fa7
TbUVI9V7aT3W4Sth4zH3FMfpnsNi5pan9GnNVNaa4JMZ73efUKBRw1CRQP2C02Z9
7bRzGdLIjimpgo8zZexKoDcD6ZDVCfwq8fnl17GxS+ysL9iKoGaxqZVRFIfxpquF
VB2IXG2+u8zpvEzvQsvXpeuOfA2HSwf2FDM0dw8/lo7zgV2I9GXhAM4umbi0BG2m
Bp7oc3Fpw4eSbuSyU0beIY3h3SFrCLqT9XuWnXX5YIhYuGZSJVfY1A2MmgsvlAH5
LC/JdszFjklCodaEZXLWKziDgXD5KPMKVFrgSs7Hx9M0dwMEnFdJTjiQFBNr4MMc
rGSHBsjT4+9b2BQA1Cmk1gg2Hy8wgI6czRKsnL9W4QrsevkNSl1+RVk4EUhWSj9G
QdZcYXMWU4GobUAzXrTgSNDapBsHZUrwnF1eIUul/gHd1D/Gw/e0spIDHSFcmjpZ
CSiDDS2OwoJwqescUCk/Upr7mch/ZKy/kEeTbvqipsMinSOEsYI1TW3HHxMvPLXN
z6F/Psrkga653orZezIeMxwstyDAhwtPsfSzUW+rspdKSR83yx8rI1L3XRbFklwB
ymP1VewMK3O3UXasZ0E0QbDqr3vNzDILQmpnvlccYIoKLPTYvFbdQU5bhTUSSWSg
XPUd4so6C7B7vCXKNe/5+gQTKJx7BFtb4Skc7yWzp37KbF2SydLPLa8w35rZJ8LB
3DPm8WKHHSdei4w2hfz/HGZeoTf7rbJysnLX1kFGuNeVQqQnx9Gr3KYxR46rBAdb
cdCAHPGVRzPOwiIj8sjeQ9ZKOUaOEx+IH8No/ndqIisn+4J+x8DgCYp1HweCNsKH
d4rRlFT5dZ7DD/AguNUwJo4nDYkVtiLimhg57uizRA8+h5xsv1ecQsNhspGlB0I8
34+f3MjiK3B58KaLA3ztnzBjg/7HCEINxiw9jap7v4UgJjsYXioSJPgkSO9y75za
ggNQSuM7RZQmkKOPzdK/Axl+yp3Nom7S9yscd0IvXhu5sgapvHIjfRkGDwjQuHSF
GOuMDlxtmI/GbnCV2kjcUY+VgIDZEoHX465NXL1W2Q9wsE0Kx1EPCPC1N2I5LlMX
zDj6XIFFaLK+Psjp5aOnkeFveadCKF3KeNiVYCWTHAnIu5QrOpEFYYqFZzBGH9go
iWpOVs5PcmJ1eQfoKdk97OMPsjFQSX8EhrEXNfTdMb4faQ6KrajBV7YZvZd7Wn7U
63ifugMZmBNfj4GHD44qYFTr5qQxBFNv9ga/3WYTRuG93skj3ckX/WoRIiM371Bj
PlzV+ZDlmNHgrRIRuAdBau9PepLT2NZaoy9zqPz311oKYlbU/k6JMjJ6SNoklKwu
/KBaIKdRPe04xTlAEaZBfMrDqu5sXAxbDIjMj2p40nAA3VUo48+Lg1MM3jZkXciX
rCNn49AH82tuCRvppOGdOagIxv0wVqIG9jp3N++TRPefkhs43VCIo7SSgIg5WIXH
2dva2w0w4D2Rlt0DcnYe+D9h4pOUTOicdIex4qieJBJU2iCjS7C2neU67NjB0Gpe
E0FL4SSstEqrATelfqxR1nEqIUg6S8V7eXuwsvqnpddhx9IrCmwrUUMYVsgbBATs
j6PKIipBrQpiLTP4Z/7mTBi4Us/tynG2ojZcM/Z1qzb7N3Bu9Fb9twVCrZthK6EN
WXov7VfqpjUzouIDKpX2qDbfw6yaDS2lxRWwfgkZ0KYoRtALCcErNuW5mN+S6OPk
mgIupTJw6l3iV7S63JOZpLIU+Kb1jakCoVPKL4RXK16YSgb9lWRTZjwAgb8PcrqN
HUmmIppPnuN4VS84bYMQjNUvfWul+WCdzLJfweaNqks0UZPxGUAgLxor4dk4TDDi
J2chfmmF1lSR9w1+xu0/Ravijsg1va8/AjoW2rTXYLMiIdWy+UUjFCJzsmE4Bbfb
3rlwwwb+1hbKKaHK/IjvGVqDCksM0tRwUMnNDBPzKYTx8PH0XWNWH7lMmkl7flF7
EJCyUZIhA0GwSRSgaFNQDAcRa1xAaYmUDSWFb4roM7hS4fPI3fYzpMynE4ZaD8VW
EO8Qmm491P4koVqaSbIjDrVmU61V2AbIETyzekvEciIwGW7MxjhGl/LYemrvduCW
vl84Qt2zgyBiRl9YLgeNJNhOFizzIY1HokEeyOlfMBHZAL2eQVltmkVwYaIDbrxp
GyNim0t3VWLd7F6BX7bMDZvc/BsIUH9jMKzoVmeY7nd5pnaj4qbkbdF80SOOBj+I
2vxdxoI9BgwWlgFEJUB8tLOv2cmhojlNJ6I1Vf2rKNzXWak6S4/obGPcwPiJ6o3S
UTf6R6kOZYYQgy8IvHB45YkM6wO+xPVkdg10omJVDdOWU5eUTwnCC8esH2EVHL9w
HTsLZ2+EG7MrVy1rgrYB/UrqvqPRdPJ9VVZB79Sf3Wf8ZIooG5LKiLwGYNAXiGhj
vMZzjQX4Op3fRw3TOMXULuNTAUcHiPNm/U2iJQ1hLftbKfokhWcQ7zJQ1/W2oyBu
zb8B/kQV1sFBeF+sYHJh8LGKhh+OH9nPf0PW7M7TSgpBmPzjefCuQZd9tfl4gN2Z
SAZgsNAkNLxEuZhABQoFbhpjkGmm1aFrjalROFu/19chIB8CKnGyJl6irDM7H98m
bZCVU+xcHWZ3iduFTffaImy2kWNVgGDwh70Rcw/fbx8Zi7Bq+pj3KKgCGphRbgY5
TyEPapDmSH+e2dBSzIcbnm8P6MyCpgIh0ib4xWDkxAfJXMvJNUYcbSUe+f03fY2n
feEldBHoWDvRaf2aWl2MZEutDIitQrEZe7uuNN2ntPhRcLYsX/GJGlg3n+SCdHsn
F8ZhzYKjzynLFwAZXzXtb7SmsGLZjMq38y+jq5X4mKRZmVG2aBSHJ33PZvKGvDRp
mDaCb8cNh0YX58ZcydMDyUl00k+ZmGPj7xK0pNnQz9H+ThXoYuTTYlFbBuB19IiF
+h0tI678d2YFOeOYMnyUBr2JxsyBv32BChVUyun+xjbo1MHg+F0EqjaQE80tGS1s
EWTKQzQx0p8TcIxnisCjC4ClwOaQWur/y3mrrAik3j4Sst22U68sSoilX0lOFF3l
4Yq9PJE60VYQbR1yBJ5hvT8t8WAnA+F/UnWkwULxdPjALHYiMIB/EJMy2yLtCVtN
Sv20dS20lNJQZ39pcjvAfCK3OOK7zCEQgZbUOUIMd+Rs2MilConWKZ9ESSSBvrGP
6ZjYsAjQdHT+YiKvbUdbxQM46OqonKBLHEAH/7FcEHK6o2z3MFwc/azyHpvCUhVa
SSYgzcFtJOElZ6LUkV9TY77ZU40d0b5s82L6650F9mm5dVDeQvURNDlxVU8filxj
ov5kgLSLmoEBQjY/GyKJMzws/SlYRLjwM48RlEqrfBSxxPz1su6alZJWDs6c+th7
wAnFcE0jax77GqHHXm4badA3uLzd7nCAXmnuuYauRDJkHxo9c0NfxXlDppf0XKaP
r4l3SjceVjkghDXG3oispqYV0DiaBGSNncjsCrN8kaP3Q78v6iWA3dRMrrJn2fet
ajmUxDYirlxtKgyHLtyXi6iFB0uJutoQLQ0nCxqqyHsKdgWsrabFr5pHlUyUbZBI
3+84fBjtVTHUMtmKnfmT0BgS1qkE3RWS2t2pQbY9DzkZ9xqn+CqLq3PYKS+tOeQX
JyezrlSDVtYyXEAElCHRgDHMQ4p9MmCZxqQIygotURq4oAF7mk6Q/Pv9WzjfogN8
cyVT01q1qZI3pdGjFKQYJVw2VOIhH5yoHxew/thWjJoO2T/BiGNSMF6TIQ/5jDkf
tpAkxzrZTAQNlBwPSIUScH90Kg9q7YRNW8I1vefPYCqDnYAflDgvY2HdgHVtIMUF
OER7/XmAo7qcxvVuej0dzyA7tEq66Kx6MANasWRO+hfhF5UuHDvxwd8kQ/islMKD
6I8xcupguXhjSSPe7YJDQxc/lESgENPOI1GRf3hONgbItJW6nQeRIKAU27d+r8mI
2U+J0MS3ZLhxDYx6HRr8/IQKWJVhyAUfJpLT1RBllNLTIRks+f250GyM05yLkPza
Bs6yN1cB5zRytU3Xl5SaICAU3F3j4seEUEqabhgaJwPdLxzOKtHtN3O7Lafj1cu/
5thfDeeSd99a75Qpxorc5jpWqrIGhy3NyARlDxTvupaRzaPNtCVL/K5t4s/ziI/O
iMN2OtjMtGdInkkTbpEXxzAW6BZSj+UvlVjyuJMxr8Mj2UYEacn+rCEAJHsGyQET
GcCKaXLxLVqkrVNsZq9il+N1XXzocaGrfB0hwI6+r9Z+ehsKpsUD0EG87HCFhHo9
7hBG3nPFRhUQCTukmbJ0i+/N1YWKdN42qRUsYDiwm5mbF0OtEGBxmszlIMNQtALB
rZ2dTTa4Fw5DWKmJqGYuNeCFxBBjGHZWrm4k+GXWM0TJbbvmRpsEXApo90TWzvky
bzkO69IaKLvYJFOZQG/MDQFJQEQnkbjP3woBoxtit7MynBFA8GWiM8VrzhMogvuY
4oSJXUpJeKy5ha9WM4c/pG6QaOHNqlilfYIbfIJmfbryLLuLoueH3vCxLsbx4hbM
bh+n3x+/yQ10iIzk84Lbmsscbs5qdoJ+kQX7ZclfVmdSk+9HhyVn2KdS/hexonfZ
ZWYvCKAn1iHFxxfC9rlQGSwcGa8OInuTGMlQuafLu5dThyumj9EuqgnO5MIswOTM
Gzq0KHtNkEREvtkguFJzJChxvvOs0EPdXmv8V/0LzGvX3delUZjv1sOy5MYlVQhz
zuH1VoU5OhjWnC4YjC4YOQJMW5cxWXTGxw48XsK+V03CJ2USV3W73EaCTzwIxUU0
AxR3siz/eYWGAan6BqM9g/U2lXp/4Ka7XjWW9PYRpPit7/m0XWmqvD+4ANkMgKwD
+1O/4XhcM+QemXcrvN5l+Mqft5TFCui28aZIsVFoEqA=
`pragma protect end_protected
