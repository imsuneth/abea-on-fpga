// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:35 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j/xU3bcu/YdGgxVydm/b2bYmJRcmeJb/sHOfh/PZWTEO8r6LdJDobqQY8wbPGfli
3UMqzxpRDsTV1E7upIz/ozzyD5fEYp5dQk4KXExJf5YI4zhz5GUhOkyI6zLqHNzy
+n4cZ9RksH4k8CeR5Kths8Bp6WVtHMFp6WzsihVjC/s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6528)
stNRPQc4w3Q5qRQohXidPBK1yv6wsOnK4dja/GxFPiiCJIcFCFUYWumaBRvjVHCo
pjTT7ThYMNTGkfSthX6Gh3IJ2NkVAyIsw2sfDZXwVTM1U6vjczqk7pqXrlxfWY1Z
RSCWHkhYtRvCBt/1E7XUKezIT1lKIoc5cWxlsp4kIPG+e0P0aWcb0gKP33q/1f4f
rcT7csF0mVKLYqTwzFVV5CEjdEcdOgHp8q2SWpCs5OXykGhpIjUg86x0EQySCXeU
0MN2siYmlEYKhurqk9zv0DJgpPkuQAT6CukwQimw9c4e4nlPZI4Dc/HUfLv5bFhL
9WWs61RyyP5tvYxcqrUExQA+8JfALUoprPqH2G92IQPAYUtW0ctQKoIdf/gT5wfn
feJRsTQxp6fJx3QH1naE8DU74bHVpLlZ84LUi1OAPWQ8xMcOG/H0Cg0a+Jtk/sAD
zWbksKV1vZ7PW8s28yr3pvFdXkQPwSkrb+VxMva9aOUvuAKrtD3H6OjcXHQDGtM8
eEBtUScbM0trIRZ4MBAYOZgWXCiDPbqmajG2sbHkXGUMGSYfEhBGEj9pO7YDW74Y
/ZTWrovOkPBEPQiW3OmpFCNJaquV3pgguRTbK+3fh7mlEJqLccBSbNI6wi+VvUij
ep/foOKcExZdWWrIhqo5qby3shNPJA5a9jTXyJQu3O42YqKnhZZRvS5GTXja1JyD
5lovk6E6TIwUNlNCe9HS/NBKgRDTGqc5G8weGJPIeNoEKvjX7t+UNvhJlTg+h83f
o0csiLHoYBaTf9bhaHZhG+L3bBAJaxRnysDxSsL/JvFSq05CXolMyyJlSrsnu5qr
ldmkBm39IcX3DBPyN0xIRna7mBGpVnstqdBCcVOZYcbQNzLJo0s6S7JJ3Kpg0k7v
TrLIbc2QL/3QI3S9vuvB4IsI+xG0SHD/cBuHpzTLSXkrGgXpOwhWnEklAPI7PIAO
ieeXZofYStKIVT1oHVDlEabVLd6HLpu5XdWfgOvBzXIqF6EDlPQ6w0izpm4uW1ag
QPd3l8InZg5sjFa0NhQRtzwJcLupgEdxSz/nIbNuV+KwmEZTatSsTus31xGPpQLX
cyvZ6uJcWs6s3I+i9rXpRdmFnLQ0cDaSccU9PqEynWZJLTUOt0kO4hmK+P8Fh9Vp
Vg5/xeJC3Ggfm6+RIPP6dDy1EVdz9mJDdReWgo786msRjmNAjIdnkTnQVvxAW0Vm
IvnMHADdZ3xdobkopI6xb0ILOBTKn8LMHdnVL89U4NBEau5oxVAjn7EwXrp6qPHC
/5sbFCGhogUbWUI/jA74RB16GN/kHOhDpyZ/v282BZvomX18m6ssHDapGn9TH+jR
ysxWls7Xv1GT2t24BM6JhPUT7U9QGgxRtiat3ApcSM4mfHYku5rUL4/uyNfwPuqc
J3OAn7JkkI3epKROnhZ7E8epGyn+sMeYnbYlPDQ+KNs68SdK0wgK6934D5d5/zno
AueN9DxVOsC3Nb+ggMG+F/u3adnUEnRO909E3W5xi/nVcKmdiqoUQJblXhMUqrEi
2s2AXQkqEJS6hYAYOnlvqm4+DFSYgNEY+HnuVYvOi305z1qgpU/glYn3D6ZO3sn+
k+TAl5pXcBG67v+AQJA8EVGHK9osq5Jal2IOEwDH2/k+mLTTaN4ZpQU6PmJyJUAl
4dnrKtN6Pcj+e8CDC8azI16rf/qTAZmfvuwY28enUlzBHJzaWmNB5QvWgOMANcWi
CXFOf+h50LFxzqYXY0cE0ed9iNx7R9+bJm6ydQdmv1ONUtHu/P/5zHJ0UUnk24cD
VVQHfVzOi9Y0Nv/ogZXyoS6T6bWeP0GmW2gXH5gLiUxsJke9JSEzgFDjul9wEgQP
WTngzz3kmjalyVScfy7DN+rIVqxdR8fwLM3niNLbFAr7VIAmb2zC6UfiJhzkmTl5
wLONMj1/XM05Um+g0UQ6J8D87KPLi/buS3tRzokgjxogjO+jnQmtVy4M6NAZCmjo
tUHZLRiG6PLmKyr26YepoE6JThhi7lrYDPn5i5eiYVtM2L7qSeQf3X7kR8L+AQAs
fm5BYdjo7pvfWRy4xJqIBs4Ynb6WnwbhUv/XhN9elROWi9ekPSQxutMl/ZH2euPC
eos5vwlHRwDR+RHOd5sihvGG6967TboETb1UbjOJMyORPRODQIMYt4+B4+UnH8s1
Q0F9FLfVFRbB42nfPXUbZZ9pbjBAQg11NeYXysedF4dR/rxwoijB33pQhp4eDnxR
/ejN3I4q2Wxz5092H7owHrJc/9rOQROszmL1auMPniYhcnT+cgUFSqMpIaNQlTxD
cHUie9VaKwltkFa1ZpcVrJsh5iuaNWdLE4Vd6XC7r6x+FLB3ne+R5H3TCLj21eZD
qr7HIBADYGV5aH7+g/W9fQ8ViWc1rAp/Phu98BqPMQfwmwXdFB9NcgR42vs//lkS
TeNTYCfx4K7+q/50wL1MH0OQL9hvSjimGX+XfyiYjymGhK0b10bqytjVp1sZxua0
wULA/qzLL2b5OOD/QdszVubsmvH4VsYibBMUxgcpaEKblzW48+dTK87pqXExrCWw
sA2tiF05tahtvq7z3CmFVyzcQq2VZRZHhXgZ3BSKaKpCETgVEY91cnJDIQi46eS/
bo9tHFxLWbkixLRS5eLEENoMgyb6lgMBmfQepnIcwfHhLN5EW2iVNLyswvM61E7A
xdCidZWu9EiNleNb8Mkw+FddeMo8a2eyUFnQcVcCYKFMsoTWM8JMzRkIE5xQSSf+
Uof1ly/oDMdVLo9vfbwH7n6uf0YDGxgg7kdWDpbBNXWRmzpOBRD+do9gD3OVpTkU
HQVRAFSAPRQ804UXS8lFYms5mfIJFkqr3C3MxesTsV/ineSKUCO2vhcRG7ssyx5H
6SnHy3QUlITSJeH+Th3mGeqEjoWWS274VXLTorMT/uIGh0wXnmPIKn23GBifcSRI
dNkKEIBf3eKbEfslK9yUnm+ylRh7szzsNTrerZpMy7VBYqrmLhbE+kmZKwtXUolk
jQXUlwaqNIucasmgWU7AcyrwzOWMzYVsHGuNLauPO8Rkk8ETVaxbH1kW8NKBs/bm
zwWqZqvptAP792DumJFN5ZKsKkf0aFMDxAEP2NkEesA/s88cCLADSk0JxoBC1BHp
b1H77niNHntQVcFvBHb9i93z+5FEJ+HB/CTrlrQ5pY4kkVBbv5MvwhtyXfzou1qt
khvU+KjCQAF6SkPoE4CqzgxjVJlwi6jrQlXyw0FqXU5qIkF9xJxsNQFmkNosDDfY
tdStSbD8Pyi1twwoTdzN40QXkyjOtks5DTWSMYl22T3kl2xHn+OpkN1rEt3cMEJo
X2eBoc3kYC1d4ve/jadvlcuPT7ufzXR/7Mb6lRQ3TEjnLV0jVlLnAZOXg1h8U74/
YfTlJkyc/SJNeE+Qe79EyEJaW/ZAYByifEgBndczlqGCKYPWYbyCNW03fP5y7XoJ
h2xasPKFLgpgFj1n0zG1te+UB1cXLHjnVESXi/3P/ttk/0BvH7VPFj8iFsBRIlW3
ZbBvrj1LlJ9lpPAvigLtRBmz4xOHJCwgfDFF84RPgd4xlh8WszU7nn4jJjz3oiMJ
o189041Ar37A8yyA4YpIapnhNgxSKFW9q/PJWqPus6+glx6GJWFWdd/7/OCu5I7C
+TSHcoQbXIfch/QwpgOXVXD5yoDiTKVO4CT/QKk/UJOo2JXBUr87rUCQ8P8ZRHAU
8K3mt5OMeLCVeD8G91wYW8aPIMjIm7eRrrOvQmKT1jFdtE0nnjr4/oSMHNxYwtHr
VjVc5c6XspPALI6dvgnMhrN4VKfY7S48Cc2uHgJvEkH4bHLnMnsrfcxjRoq/SnbK
dOjTurgFR8KEBxGpU8nJGn8GJSV9pRFoeMJoOdM++Mo64n4M4WyIb5u9fhl5594z
IWksCFZbT7dMctr53inN4wS0H/zMsxRG4GS9mI3h9Xt+M8bGHbZGtjqmhCptzxyR
8sh6OLC8QYV7HT2+0xRbHc7YRDyO1I0eENhbX7YWQ1cCHenp2h7OQbE8sPdtd4/q
Sr3Mls1rB13AzTjJNo8CRKA9aiC84NnnjpzHtGbC8kPlGh0ces9OZ7khl8taV/n2
cIfisJtghWilySws3Wr+3iFFpqXRhhvKmZ0jjyW1zLdBSj8O6TAhmwNoYrmZciBf
KhAeA6RJMuLQG7o9q5Motz5Xd0SacrRXqnxylmlzPZ7jfi4SIACJewfzaNCvinnr
GSWu9sFK0cvbNBBx0ax4FZjsHlQHAelHhuMHlN6kQ6RR3WAAVuw99in/1fQK7Uc8
ea96B6MNjRqf8C3Jy7j7TZyW0EqgceDIifO7FDCX8xbS9kavgbsxPcYCtR0OARCL
imbMcr8IGAR/ut+bTxWzuqZSv7I8JA5YV/LwdX0Sjj12jHKodXEsXliwx+Ttvmlf
Z1tm9uoRUDSkuvJsU/y2n+eBJ/4OOgjfbaRTjrdRoj5yOFVKcZHJgWRixed4gTNf
dOmRkY7ILhFGG9pFWiQYJsfHFTsJHYoUtmZmdM8Kc+EIRr1+201lDvIpasq7yJef
bkWu9L6oot8VOILS1Ymi7Zv+bqaMzxWj27doI4SkQISaDE2Yxw9ZnbqtvdjmOkw0
C36XoIrguzbKmlVg54k/rMrbiQKlXi88b5NkeM3OWtLOPMd6KB3jzLej3QsLfxXO
6aVWaWpp2CR0izAQOp9+gp0DS+Imw37GItvJBpLMy/CpPuB5C486Pz2zI6MNN5IC
bQcQcyWLUqlm2HLeSvMBSmAXUO6QBBD3hZ6f/TmxyWRVxh11yhO4DExccqUcA7tp
asvM2/Igf2Zgv6ZKupjuFWzxjyA8ssL2iftia0k6dtnlr8eZC67q0EFFYZn8kauV
Df62g9EFQirFyfq7r4vCqgukScuMCeSWJ90oGVTyFoaKUi/eGsnPhcCpd7QL29c8
qdMOf+iGICyQycFAYzo5HdMAAATApB/LjlOWlOTe4ATZySCfEl5K4al8CkD82d82
Bg47LRlqksJjpwOy3JJSv0MTSUlN+9r2IbGne0uSdRHQZcOtsdTzLFBQ/AfoI5Mc
7mJor2qh0g/2oiMDrW4js1OXKkZsQFhE2/gDLeuAbLipHiTtLheRUH6qyaeV3Cfu
NjE73xnziOPB5OmlEjM/zMO1e3HjVDD7pMRulv9M7kAdvRLgZIYgJ3t2bH+T0PKC
F7TCgpmnNCrRmXuoEGHQGfNgVDjKgJDl9FfKOHmQoc5NyN1PANE0+iensAIPj06E
a78rlIvGqnVmqFdjJRB0bxVUV6N8JWnn7tFRNTPkrZz5EX8Z18/E2UFlkz8hp95M
332bBqeA3qY3byOh/c9k+QbdM5DWiGp5paw7z01DnkeL46g4elgs0LmCXTAYXJcu
25aBbHG+LmvIB9EXFLNAkocJzEktOjflc9j+32/mikNzJ5mQEzWEGHPzX1/1sjb7
acMwFAcUvdxwTn9E1DfC2DRZh5UYwkVF+fJbZSPMY/+pzdjo7aSA2R24JmJBRWmh
fMh/Mbg7wnYjPA+o//Oy8GsGQ3zEF209C+UT2RZq938YCJUWLV6rxXppon3PdG7h
yjPd0ynAJMSiWBoLtyRAGBYjLnNjhjBKXy8Fro/REWUGMKfovT3A9H/+ZLDhvSn2
WdI/uXMcn6S7ZvW9hT4YXMCKUiTPP5C71WNbn50hZTRslVF8vNYRdwPx4uZQmBVS
FJX4OYG5gF8TestM6ESXDmLgJJoWyj9ItstI+/XXGrBKZgiUtYi+EqyZB1Lqf8wl
XeC20KeMmqAzCweBvl6WXz70QGpTldQLEk+N4OXty3F9pI40S9kyZJVGxGPUCffn
iY/5xoU232GyogzwL0kkhiNm/BXcV0/S2IF6pbnPKf9Xfzozm8QRboC3AOjHgmcn
tFPO2TZ75Uj/tubDc7u6T629+n8aWPyU80nli1K8cdfkC9NyJwqyKmOdzOuVJ1j2
2aELgvn8yIeHvzTZghgU49FoDhi+pGKB3r3DtJT7Ll/Ue8pKUtknFO6JLwsY3PA2
Z58NN93QI3RWfhVgZEztte0SPED+sxCmefBEQKZVXL6e1RIOV5LYdDu9Ag+ZvdDX
8C9bFSg+CPPHAPZetqa64CdAJrn0A5I/NquXpLz0TEx97cufPXSrxN1+QXoqQb3i
OIobYlq5L/oJ/ByhAdch8W/JHcr5HvQeE7q7WGHGUwmkhnUWzBp1nPWGzV1ZQk/L
awC26p/YgHlUe1vjnJtmWp2m3y61mM+riWGHidvjbeluAxgoO43vI2fPxOr6JMfO
GdcS1RBX7+V4v2gAIqYgrpyknkx/8sou53HyHk4+6fjYK0Ul0vuC/M0mp99mKev0
5G8iPb40Ml6D2HaHDd0Dx9n6AkwHzBQE3wxNqIUpkExJUsuf4VTkfIehmpt8RiEg
ikqcRn+NbThJ+V5jCVsXnf4E+1xaLquK5ECUtnEfL4xNSQI4YIrFzOGrQO0sNe6o
aC/I558cbyhcGYMdV3CZOCkY2rQCfFICBNfdzzG1qvZ7svizu+7gtuo4oJOtLyR1
9LiyiqKgQpBxNBFX0zKYPzM0bDIuptcrOEGy0tkVjVTQvBrIz/tp869nYblbfJde
ttNJZZUWKum2RRGvd3g09fudnX/GIUibCPW39hNxNWFEWdy56Qcc4YrRo5O031Vz
WfPvN8zD9uTgENJJEZBf1su81ULx13nvUNVBzZjsvMdGkv4ZUXj+HdLT9mxwmT9w
cmX+fJGZiGkfHjwJAX3wfV/ITVul2t1OqDurQ0TxjhSmBxK+KkylkmBO3bqXnVyZ
z5vSZrCaAZl9CZKqn/wcqfe18ixBDUCUzlFLzR8mHWvqXpHrwsZ+w+pRIvzENOnh
fnC+Sp40C7FwAI8653s+RVZfAKHw2poSKN1ZqdL6rPIxAxK63JlgGFxW62lVBKZT
ishZ+M4b73UJ2pV78sFrlux79dqFO3VIFjQxtlAlvGQDEnLIOBFxUPT59av6ECp+
6mnZ+zMG2bCbVK9LkB/oLtbQKxo5yft3/yeITdDRCu2B/7uk0RbiqK4xIgukXUk4
zlOcMCt0JaO3429jE0IaShPT+/cF9nwKINokJKKzSW4ZyVszI9AbRDGAq4cJR3rU
ScS3hhVbpXNJ0qdgLqpNNAImVfxv1Q8Xrvm8JFD3iq8NTC51Hyh2ROr6dzXQrj70
NB6yUuTwLA/fcUV1NCDWl46MexIWoaFSZKR9pUbn1hTdn0XFGEF1wbQyy78X6rTV
PQw9iNhuLl+SX/f43qw2UodXjxGfkRqZQOEWKj9vm+NPuMeXYqIrXNV4E7/FsaA7
Wgus+dE/zqJVOuETCwtYYOZ11Xi7QPqwdXqD32haTkMILCgjytIIvTp01IrmoyUi
1rvY+5q3OdnHd65mGalO2dVgsQlGhGfRcH8P8m2yTBOBb+axjlv6rbXWROw3AGnr
BxTvgCKeFLW/LgufueDk5clxEiSTgpjb+G7Im9FfjSLYTOEQhvZX8uSpvNiqcL0x
OxFnWsOnPkA3Lvxx5rHoliHJAl/ybx4tyYJEITWyROoNWx/ZzGAldGQAyvTDAxz4
BLLwem5NhiHV3OTQYg1LizOtjf4hmXmuILShG1xuS4CW70x+pj67mSosOxVYljiK
PBCD/NZ0N/OZw7+264Y3++hxS2YDqMOGdo1//hgs5uGGHwxTRYFg1rBDFtVyeFro
93G9J95PLRvOEJ1bKDYtuMRj33SNIYQSGveWAVBYJ3VnsLMUMBjXFXj7/13eQ4eU
Yuqa/wxl651pv8QH9PhaJJyVhmzzUmnCb4xdBEtA+FlhC2kCv4vxWFMD4NkoTeLa
cqMf9QUgzmXxLnnX5GooLZHv7jQKuEQhn+MSKRar88HsT29fNqJIaWohQXfAnWOo
0MQQAx1fhzSVkSVeDMZEJOjD6VY/t3c6obBXH7RCObDAB251CdhtA6jGzWepEwkd
GttEtaJv2DSSnHOgOUWu+Mryyf+SDJPWlhiYpW0IA3sLfD+PvR3KQveh33wAlprB
27g2GhVWdTFXXEnrat7ksM5IHq8hSveXvwIyLXsfApsYM4lj+MDeTJLXV9lz7SJw
erLRZ/45XGjCybzAX8XR7//tbCOalTDZ5bBD0vkIw0VAnxEJcM4JycrMIET/dcfs
R/y4oCALSj9Y6t/greJO2GhThxOBseGDyGt/6eEG1yt6tu1XfGnXLNPfsQXuo4M8
5EEEF6M4QS+hrq6IKCwxyC1e4g7VIBaPPYXBZEr8AFCCxn3XD4fBnsdpfGApMeex
P8wt2QNkqYywlErKB+InOp+FSiVM7V0hQITuSoqR6eW+gTEswoweEJDIYFGCpd+A
aTqxKc+mMUq134AK27Fk2/4zk6q9KoGOfICuWzXXVcrO/oJZ7ej6ozuenBQ4KsT6
K4U9xlPSljIWwNQKxbkTPV42hK2LS4nN5ipvZnqym/Kpe/uKYsIarzj9BHFLgS8V
hFM2/nCXJD1mc6oX31nYTKxcLM0bhfzMqyldn08gsApkPj1BAUyg3AzrJMNwap6B
LhpJsr9LKe3eobg35cnrflyVu9+ZoZ6Wu0pUEZ1CSSoaWXYxObza91/fVomBFLVU
wETotye7IJyWWSET2qqqHgePvWbDJ7xX8ywIhSOCwzHo1iqDpREQWoRE2ci8nQ5d
Un+PxU+fbwuYFCHvqrS4Z04FwUcnf4fkkBqwdqawZHk6P8zM8uL+NJmBtVYPoxQb
`pragma protect end_protected
