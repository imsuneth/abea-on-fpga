// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:42 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G/vjq5ZsX89GR35ARRfP85XFEiqZdkeYyHmcSsNfMGpHFXrvkNvV1M6pYGk6dtjR
8L9F0Nb6v1fJxorq4Sb38ARhTB7oZ5voahz6o/Lu2h/CH3ig9CXgAe4HngyEDB/D
5EeoNWi3J9WxbJ+DXLMAJqAx1zy+NgYicGmqWNU5oD4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11296)
UZGXBvakgI+CaVEHOkAmPosBgsM0Gft9k2alKTFK7xvwnqb74ruoRi+UGtAooUUi
LLQxcmSc+dQJmqarArTTAWoNHY47v1+Yys6YSiN28xH28VHEWhcdqeUR78i5epvN
3IKaURCbYVtsEwPQMIgcUgHOChXqnDbCSaMxdqX/vvcH+Ximhv7DOPONOf1Zt6K5
Pt03d0uMAiiAfWug//E07zykShQFvdp1H7oIuhzWjhqs3l9ZGd6dtlFDoLH9fhxz
J3wvZgtJ5uhJicaR8jSKz33pOsa4zBO95uw35XafTBI4BKHW8slMrOs+zYjq9N+h
J+BpE3mlfmHne02dPy6Dv0QIgS72w0tP6WuF6uJ+BcBpPHudTgjHsY5O4FwBmPZC
rAcxXL1cUx5B50nVYvp6ccko8MQ74L6TpnCVu76QMzExQ58VW/kmOuXpgvZRKPFl
bt7kgI1XMhP8K2QTqUXl8v4qhDdQch3McMnERPPKxl6v8xfoH/MCS6S4F+LtGQxk
c+fGVOrHvmY4oqW1Bhd9T5c055IITreS5a8UrFfvd73xAqzvlrY7vrg/hac/1m70
G2/4gwMth4D9B6MiMmGayoVNMo064dd8OpRFL3vL/8t5/ixxQ8+KpyaPEfeABsWF
ZqVumpyzoDLoo0iDK7sBPbZ3qR9g18GuNw7Y1DD88fPdJUJb4ixoby7/KbHXn72E
YwCWIqo2OzhZ0SOufmhGaJJQ6bgmrVJHn0/Q2VnHzC3GckwQ2u5YeMkm/althMEa
GplKotTWxSZ3HD9rJvdtf8QlNFC+WnaoZhNJPkWc4g/aYObPvkcUzpqyKnZnoHD6
d+4rw2zu8r0zZG7MbV27Nyt3LT+BFE3awo+D041S7/I2CPe8QODrkrTYds4KnjAC
Arljyqe9v/XcGCwHQHjJDvGVzfg0c9VuIKRjkVMQr0L4Dn181ziMWA1chcItvcAA
W8Oh5Z2x8JuhNkJYXduP5EcYgkm0PmIRXsl7Ru/k7tEJ/zdYKL/Jti2ElF7IWq3F
f3t7MZkfrOXiz9KNefCWN648LbDXxUpYr+00Jk2h4u0gWezAzwVGzYbVWkrx12+G
qIYDfvE8nTUBw/gA+ztROzoEBjafZulFXqjZvNBOEtQoGgzv2tzkxaZyHHL2K6wO
G2RQq8ePljhu5eOnZFbYSXBXCP499jbgOvvQiv3wZipQkn5yxVKitEtDE9wgMpTK
ODcwQg67r3oK34WP3ytGlumXm0RN+1fDBbVIFTPoAEb+fiNagP5K4C/yrc6PAAiH
3yD6KMuChl7rpnxpMabBBSIfcuw+A5dpZBJM4YJpXHvMPpbyTB7pLD+yumMNuLMz
G3Qqntn1v6iO0EzEmLZ/dYpXE65QSeBCCzf1BBuF4RPcMYz3lRXyKkWop8JvWD2S
kqcbl/1d+vr275ODXB7X2x128jmOAXDgusRzHNy0SRrAcLtoDx++quPDngUGe9j+
HOI4rXkdupJvNrJ0ktoqReSWvz+eSZl7CTOncadd2LPg33NVgVUKKOHwaKONUHCA
1eZ4DRKonzcRDSiuXZbKAlqr6E/wf+tPvoXhs/FKAoaLa0NKdN0MSQ6vjGI7t1Xx
lmR7y5zFDtC7kdsi/oFXWuKVV85FYwOjKqlBOrT5h2PkLGeaLwKHMFDKmq6D7CDB
r273NAnpwvCl8vc6ZbNNPoIWWD3cMyx/3nB9htmpepwxhQiEtp/eTc8LqHXc/TUq
pM/gJJhzPb7y/8t+0LKJ5Y9b4pahwZslvZ8AtbTP2vDZ5AsYlYLrPvLCL9lxkLrv
bbp/9zGZ3M3Nh/Ugp5z6rFrinMB0BcTvs13OaM2HpRVxOoUQlrJN1uN2jL7gJ5NC
H3UGxJ8ZKRWDgchjKBQrIieD25I4frsSpWQ+ixtm29LCceb5n67uRCTN/CVYEq1H
+jY8LWOk3CXUadqiVVTZxar82XREvTctHZzqT/4TLPJ4xeBfUU84nhDRBhfoa7W1
F6CP/6a7v7+RTmJghLw+Pqm4wEUoRT2e6gcT5xdP0SjXo8ptoPLVgj0MaYkETnmC
oLVEzZ4w4M50bUWqZ6OjSNXU0UJp5/dWrRtwpYzk80pXzC2u2lnJXIS8pZUPcOpq
BQ0EdSItmDmATKxVHx/nUD80QyzcvRSwEWdNBOWJeGnvrejeH8e3i234dttsNWXo
I4UcMgunVSx5MNl7+t1plIvEfc0GSsPdf1cc8mcVTRAVQGSBHDbS5bFiQvCyRnFy
uV6N6yMZgaEnU+BsQNFiftPUhT4AC/ai5KnnB6gsJq6wZfAMrtH8a31mGl49VDHy
tcT5uDgKOfFuHqgSgJwU49s9J3HExYQ+fPUh96rJ5pLrFJTAZBIg67pLMYuX7+jY
qfRznpGqnGlxc4lddDIlACa5OIyA+uCwaycywfBnV7EsvviZPBWBPlqtplcwLGPQ
zCt49nzzC3QkLu8vxuecdR5vwFHO7VhDscoYOVnDgEhVAYEo8iIIEgjMu+vWYgnA
8Nd3CXU6bx4yU4KNaN9uC800pIBLx8oE50lGYATulrqeB/C+L52kexcxTe3AeLYq
fRHUen9A+HVNQ/6R3mAK8uA9sYqqCDrqyn4OEyL8/mDH64ZqESST+BAoMoHyoNhJ
9zdYgHE495T7lMmeAjZsbZRyFEIslFTqmFH8BF2XVyaeZa7eNhaV2yR515y1Z4rs
UaUf5C2Y6mR68nFPz6K9/lJ/a2ONo+fMzoEWbxElW7+4a0RelZbo0SbWtTW0vEFr
2mAhcoGYG/OS6Bq1QG0gCQ7XdkAGPzG5IjNlxFGkMkVa88xo8HFYN5qDKUVLupPJ
SSqLfr63HfWbXZf43vqsbsPsPiU/gELXHDbdk5c0Ug7bFWMPAzzxfH6nuEUkCrkn
UWm6Cqurxk7jtE3jli0R50BlBNpiv3yMcyoEuBDthYo3NHIrYC1mvNnJOpF3+UzT
eADOrxYI6rk7kR3URqAdQBh3dt+rZG5+TKYb+W3krCHncCBYRWlGPxOVNBPmGchw
9SsDuDMun1h3FNkCuUy7S5PwiMwiqLdp4nfzz+33n76T4gcYIaXOCN/Jy74AmZFx
ZnFDPRcLpnSDNhTzA8lPstoYhbkF0VRbg599I1dpdCvfxYZ0lb4JpvIBs6JfP3HL
8kJrfM+Mo5xAbDiloWT16mx3tV1Qc4zPS+sFXTtO+vXFzbDQ+A13GjS9Fvy3ugiz
KRT31VMYpkNHfaq1Fyc1aDAPYVN/ruDUZmSovm8T2RabaJdMUDoOkPYAOjUjBAH+
DpjZu7LRe/zEvtcATbtN4CNWMbTwmuUHGE1NvE1XSiGbcUjX8SF0OjmHEv3iBbmi
24mSdAL3atKoLaURFHdQwyq4+ajnFx4dJrlp1hrWWVatySU5Luk3+jXO8aMPiiVC
9hBaTPVaYsm0XuDA3vR+hNkqB17SRsE1jwU2JGxgWlXwVDAMLqkcNW9fIe2H7onj
rvG8dqHbZpkQVb0o9KjP4zNbnxo1X4dBB3mL5afepUkI1ow0aCHT9qBVwkrAt0MB
zDwZ3CuH1R53EcN8e/u39wJuT7LsSXcOoBeY8yY9xtV7ce9SJIuDaUPvUzyh1Q4A
n/q+JQQycIc+XlPPa5c2azwAoSQoNW+3/Q4ojMYcirI6JYLlihiVksSf0yQOZnB+
6Bu9MBwKXET7hmT5KJtrrIIOus+J4dBWJzx49VXhwM386HwxNqRwM5tIXIJcyjLE
JWMeQDj9FeWi7GoEmU6lUMP/oDwj9Jh7hJv6d0htZiVN7YZmROSWurHi0Pm7sVx2
3D5s0qZ1Hx1fIicZ6VwTlUcLX4lbnZ4HgposQrTvlbAoCkeNUjnKJAUNXbEKB8bR
KxIljI+N7DkCFece5ox0YY9f9Ct9ehcqY6Ltet2rBx+MjfHIV7Ta49grJl1XaM3u
fKf3mlwowqrfI8Lgft5r0aHFXJ/pfVhvUNsu84u9p2/diEq/i8qy0FR3+UtZq9oE
XUrJ2pQptbs8xRXZ4ulK9Dox6nNY+b/04qj2nZgnK2fTzc8Yoad/U5gFrAp76g83
PD6cm5BUmxdjDlSS/Gs0a6+Z7rDJen0OBZN5trc2TMLgee4AtrZXq0wMC1TLXSne
iuDs8REkZArn9t1XEy8frnfDYXq3JdyiXt4BisDxz4w/Zp7VZPkEtU/6Lro8pFn4
SEAg9l8JMKZ9XvZGY03utXJ7Wg4eEthJZfBjgtOqBWrd15NwSe93VR61SGoozsn+
zkYB0f8FvULGDnTUNdD3DrDK+Zqrt7SP8r2s9OvLhE5DVdgrOJClKV+N0D9yRPQB
N7783SKXl00ytVuiRmb/tIgCGrXz+BsB95wWEPhnZhntmtHqMa6NFNyGLXqWhRPG
n3Btq45X8ModjvK/VF7mDp35+EIjvR2QiLsHzlRyR/T+UTvjknsbBJLEKKh0JIhn
s9tZ/FPIzmfliuWrtCc8ayR6B5Pjo2rsO4sg5w/KhykvKvalkP5gDXAKdxQ0EfFZ
LsalXq8c/fWrsgLhsFFUzlqlzSNY7WYGH6umLhGJNFM4RvvU7rtsfpyF3blYaXlg
m6b5DP2h5TCVFnrCKDDR/RnkF0ZV1ps9pUrvnvrCG1g4UfbKcClIrVlkDxXSDJQO
EPekHEEBaF4ngHgMuwORp8fvb/44eYj/d4F6o0n1J3IEeD5thkTPp6vBmmrAeuqu
NJCpL1depY3FPrqw2ADjlWgvDCEq9hB7cLpD31MrUs+fACFhtaxIQa2HcIs6/cn7
oWwiSILyhHJrsBABHKXv3lTa0m2iyY7YHIFuYLQOU1o8TmM0w0SkFpzo45MNF8uo
W+m2AuaZEBEt9qN5qlDlkCAptmfWXCr/agiFm4ebeYY8UZ8eB/shJa/fzNFeRcoq
h7IaE92PbAwR1TcoQ2XPU93pPe9C8cOyzRLngFvsqFoBmd9fhJK4FrNqYGxLJM9C
UpwQYT7hJCujIh63HhXdYeaRoxmKURh0XJY0Wk0XeXg5z6914JHI6AeLZkolEb8m
KQPADwpoqLqgvtolHq18yJUsMskFd85Oc4NNex7bKNWbi9SjS45Pbo0nYzfVDS4n
TWn9m/VuW879DKkMzdMEZJ4arXKg2+rXDPbeJLuqcHJERz85Q1gjRAoOmwlwaCuv
eEsaWw83aypUehZc5KliEuQtG4RUB4Pa63YPLMXkpEKMqxsnqdwGu6zzKlU77Omc
RamvP8yc+8qCJvuLICoW+9op3TPNss4u+lb7gr/3mBtzMoi0HAKSuIV1PSSy/sWq
St0fgByql6/sY41WzGqakEYxq/vNvgwTK/BSlC2lZceWQkFXZYiu6iz7A7ygxU29
iNgPNNyGIUZ2EmxMP3Ty6lAUMKlrhhLtrmgOUkZBm+nNb0isN0lFWoKTLfG5WEnu
xpdkAl05bClC+DqZHFHeW+Xbxz2c4uanTpqMjppp2iM6a2iYD/yRirBemlv/KnFV
8aIRE1cPIWciClqjNz5uWbQ1Jb9i3i3JC4E1G7g/PUCy7fBWYnqjijzADU/qePrQ
7awILtu0ek6WnnZ+ez5RXTw9Rxf/Q+BfltpSdR6jzDVwZyMqoUPypkuBrKiEmYq7
b9Msp5HmSBnAauHZTn+Am4ogIphV/NgNOEEEsUM2Hp/q2DSCzvJYdiWAiVtQTTif
0dS+G6YJ2t9GrULWfcYjkgDe9sIQLB3rAFtag7w98A0skaDGG2Q2Mo2oary1OSjT
Taa4OQzRJiptusS7G859NKN9dzn+yTgcYDsV8xHzNHie3V+pLTF3mQ9vNxNCKdn5
9GI0ldCC9Ccerx5d7+AN470c9vONQ6pmfMILAgKKS+tRS+1vb139OGlg7fHjlYuH
UhU8Ixh7VmDjgSV/czVJ07aPXG0ONSfT7++AMH6HKAn2dpshhg1Geo8r4D014ccF
bzEHZF0gF6uqIXgkfeP/PVM8apXHBaNgbsc1Yf9KGmhXc5JU0Ym4n+LljE9jCszt
PGirouIo85GpDtcymamGXGm4U4HwcvBxJ4Wk+pQ5L4pnSt32kPgfv3n/IE/y9ZF7
Cn7fPNv08SBYtGX9kPw/Mk0Mtdmm02sWhjf8USXTQXQaJXt9Qok3P6QWG2z8rZSP
3kvSZosWowQZ3KI576aG+nVcOm4Ru+gqRPYsGGBJ4+D4sk6vDAfsTujZjL6pF0LP
Req3Sc80bzMcZyRVHs6WWhDRSEpYajLe8tpIkETie5Xhr7FcjlEAl0Cz14Xj5sEz
M0N4rHWcEAn9C7r+YlyOeAqIaD7F+pnPyBu77ksfy7nzHl+6H8o/k4a4EquwK6Em
pYPLBwHfgc+AHcihDydaETsM8GF6NyBx55b+eIeVmcYrXLbfaGrt1w9sQlVA9wh1
oig39xYTVSeDqA79GjasHBt4f2lnwZb97wkvHjnG60bhNidb7SeVk39rP6V3DqNn
2nkU6tAH6/dAq8X7svRXwVUq5iWK74QAozSb1wEoQkm2attzWyUA8zQ+GR4ND6Eo
iNE4NAoow12GBazcXKK03qdj6w79d3oQw0JrlxDU2Kg9+M3XBEWK663HkKXp/RGl
H34NATtOKBCSr1ar4WyTr/4+V7/+YaJoHNDWjyj6zzj6hD6JGynjQZRgVbNT9/hR
HmDN/igKYdR7UskaoiuIaCXQvBdPvGaU3mFKpMMGbuXFEvz24bLkWGyWLgX1xyMX
h47iD5kV/pnkZYi1GZ9b6CMHZXDSh0asWQP/ParRgG3MGYBkGWaSuN82d6i5A7TP
TXAP+aWD6rX47MepdD8d3vmMXmRTdLnTveiZQ+qIQxOFBkshvg1+ML5pbpE8hbvS
cOjEo5jEcVEP4pRcUjxD7+uFSaZ55WnTNHoiIyCZgDEyKRbaykdd59lWMSW3MCfE
jHceGPMEbLKyX0LFzyICzQ2y6/hpN3+C3u+BGwCkMbYJ8IzfG+r+Rfc6bprtP7wk
AHfLqGb+mLy4p5ovLP9rtB0bBxpAYQBXCOKEhv4t+tc12szOAhbwPDZ4bcmdxTxl
HWezb/WiNOmPwlA8vj4EjNcN9hqc3rXWZBqsC6ASvxzd9mPUvTam480W517Rxsvo
W7jxQ1e4sD+jtI0F4v4XaweJ2Ct3xJMqg1LIyxlGAbxSLghFTeWTpMjcBQ/s838M
AywEwBG6TLRD6kiXReNGRW65pQz4DM2fZ0iyVePPcXUALtxlnqtvuPaD44Or+eac
6nal/0S3ry0GtuIAoWkciwLUZ/FzLjVtJeEKxcuRdlWoMKqRaSgzjIQfDa/oi0V0
EXDNO7JlDhbWTBZcVnb1JdmmQegd3MORYT7kFk5gD9SolIaQuOR4RYr1bt+Ghfcq
fEHXA+KrCanGmG/7o/Z72r6XVGPe8A9dKNCv9lN84/5wTS+vKzzEUTkaf2NLR978
IFRkkcgbC/wNMY+IWbbp7im932e+keGoSPbaCxzjkh6opPHmSbVtBDX7Do6uZD66
xYMldbPI7J+ZfH9GrFXkh+R/iyuDVJCdiBqOtGp/eigoeEQp5ABv/RvVCEpj6BA4
4bsxLFwLuksuNgYWZdPy2/sB2PJFUtLxw4Y+rVm9ed0gvzIoWVwUljnUHBQ6pFiV
ODrwK8rne6DBj4xydkbvTmWAgcozIs/zrTidX1xzSaLPsisUc1ZL3Eo94L6gmetE
mpjbOjuyvM5mGaKHj3ou+t+S9/hnih3ReNygA10XTj4PcRLdkhPgUHyYF9hLe06D
HKLOOD3B6qN59V8dP7b9nLSUx/mC4oGrefZL+ZZ4ncjopBon6Gf3K8ckh8vym6dL
O8Ike42sX/7zGI5inDO20SfEllwk7JKeRb947++/rJonKOv68O6rxnjNjLRyYZhf
xzxIm5jJv7poVWW0F0IUi1ckd7Psm9Me1noh0TmyG7wVfGf9UjDZhQR6JeudWHEK
OKwjhWtdt1PBu4t9tgGCwLp2GM5/lmXr3CpfSxaNsoUOFVOajljhiy5K4oFj9uQc
lbxhDiFK7DwrgkLgOCZv5dK1fxb/WanuNwS9b//xTSgOeDmPV836UYDgHSczDLDH
hov+BAN0QOq62AiCe0kJShf4GegknhZmrS73RAW9C8wy+xeiJSkTM69qvsnLsJeT
VpTx/NCWkxPkPwGew87lE9Lga6nM1t/uxsK6J/gf/0F51YxnP+7PfabkHd/uh6Mk
eUmizNBA8oM3hk2rel42NNty+W+uMYq9rIUtTFP7z6SBerNmpGAvm/csCzi3ihSg
74XMvnj3xN5/lsXH54Ym8RXYX0Tc48iLkNWEP0RSlL4Y0BFeOFnH8dUc1vvlQrWM
Q9qGOtzDRjGmv6eTofNU8ezEmV4lBKmr87gwGVOpuhnhKO6WkUTYm2ymm3m2A/Dy
RePTe+8hzYY1C/7OBq2lL7yqHBIqQEBR6c39S7A3qeaCLE4WOEH8QIRcNqLB6v4Z
6bo/MIQuMN2TRTPD9Kr/SgMaN4ALFo9HP0QF+RrUoHpHJa1heT113g6sEo01oiDt
WfSnlK8a6bX5aeD7NfA89H+wbxGCFiyxegdsplobuuyzg0lXPeJRWm7ILR0cl+aO
n9dhRMSUZlG/WsCOGC4bZQoWqhZzbv7sPR0sSZhxgFcL+rwUdRuHElX4vRxw/i9m
nr0D0GN3AL8/P4FMnhB9EpJCJchlFVvVCw8nKSL29y3NzZJV1tI0AYMAI1p2OEfI
mVRTTgU/X52VHar1aSzBLcaqQhhlSOLbLX14h8uDmRXN97zHcmYSP7Cf+3i0zsbK
ygaho8HOhrBQL24o39GiRCp9c2l1JJabyN44oWv7nEq1CQHcAOlSjC3elOV4W4jr
SfCXe4SCa8lHqwHoh1VseHpeuIaZ5nhYGQ4R37p/YMKxNfOEmsHcw36/sRtbApcy
qt/wR0Bwp9yJMSqydOo83RcmYeZZ+HD9iXEBucv4SBVlJ5pUC+rSB9fiAe7an7nA
HO2dFQpArNsb7VfXkS2LHPIog9ijYkFvlBWeb3qm4EkI0wWfM+P5R/a4Flqbq7B9
1ZkF+pJSG1KHeGv21F8N+T1pBrDnQkfhK6NRGV5qda0VD3fhh9RkVOk8bhzE+KMV
L+675P0/M39QweiHJV+h2rARvyp8gnhZUT9H//8OKyxVVZaia/R0N/0MJIiSOppG
FO2mN193EE4byO023ioo15AyWWFq82fBeg6zCJilnosDWfqoZB/AP/XVIIhGprUk
o40Dr/teGixRlsaXE84x7Qu/Hf/jeuGH+9xj9a4ayCoFVT3xge9fpiZ0yXJsYSc5
Xmqd0jCGPGsk+YQdr1n5YqKPRASf8aruEBLoZqBtcck0XeJ+O+5C6e895CiAnFf2
nyub94SGWpUh9jIQe49e3oF7shWggwy389A4CtGn6SbmR1KJKWs+SesP7M1t3j4l
y4YXVXj/7OuqMeGJmbpQ6VYY3BNS+o3jpAccXOEAv+pzLluDeArX8CyTwn1TGtH/
hxAcGHp53NwDIRBodGMdfDDebZGvb3qe7XExP8hqagLNhdosknxIUrq1Y+ipgQlw
drNU1iubWP7oRLR3lCMu6zCsbBKA4MmCnXyh7pk8witIXcHqA3Vgs4fN+9KTgacW
D4vqRVt/ByUNnWKS/PgRwGGb8K+vkaFZ7JChUImITDHOA8CiS3vsrY8xZbt1Nefa
m/CDVlijjJzjbUDf+Ss/9sPAN01ge0ediVHJX2FuscNbe520xyy+6iuDT4w6GL03
S/cNynCim2GQT9kZamGqXSA7v32LFJxl6TlaFexrb5V96vwOsj0X+5PJlxKYcsFZ
LuPKXSF5jyXsOHBhzYhCjIW6RXFfj8JVbBVWxxc7WZ4I/PdvuPE8dYONf8UzHkTE
KoNi2WomIpIHLD8zHVjVj1K9/0aTE8cX3f5bNBJbFKhS5Hf1tKfn2Ya7NKZ+bKli
66FYW/62em544o+YYyyQuICWyvs3gL2wrwpO8a2+wanZ0taV0iJ8G5otwXCGNLyZ
28xlDsg2e1pA66ZpJ3UVyWuImtfcEa3ebdg2bm+bN8PVFjBllJXtEjAxL8h3Bp/n
sBRr3zGfXS9msRfU/tYxrqYYNlnvAmsv8ItX/NydSxBK998T8tR58DwnY0mp3Jm9
D0eU0zb8D0NfANruWUvdD5spLQWbSdv64/m6ndn94oN0qRI9pWXkrJ8Vo5yneeiq
ldMUY4ZP0vpGKlhC1X7WqwUv4hd2aQlDHFsq2y5RqvVcpZOtESkOpnAF7uUSaOfm
y4gkx6hB08pQhjKzpIQYB5MODKllLuek/CRfUQpynFIIAo5FPaIQw5JAJVWWgulE
qRERR4gkG3DuIIK7M6TBnEIxdGb90g3GT2q+/wwcfTPaKfFqzaiHCsrW22Ssahd/
2D2K0ghUHIJBX5OidfaY4N5o7e4RYDQsMaOR7f9QbXeFkDJXaebmUv9A7NTr0Nfl
w2xdiCC2+XS8GoTXn2e4PVzqTL0AhKRwlWIAvE2H2LIu6sgNOXmT1uCMabSfSa3D
fu4vCBqZhtb/TptRTjYxkVeJmfLD0QE1SCK6PBhvIxIBQCjpzqDOYFrr8PzKtHds
ZHWX9QfKXJZTA2TXVe9uDpU5IpLMk2qcjfRbyGDlWhVVgEvc5cBVYaTBwSq/klQ7
X7Y2bQ+lqHOtrRRSIcPrwE/e8YS7FN4a4bfkcvBz6+JesvAg1Sb0+7AjGwbrgmKl
rBgIc6GEfC2uUfkojx6TJvkeWpqPBeJKJB880OSHXJPLt7vMxJc2+/8blFaAfttX
g7S0L6cgmgyGHXeyoEPlYxdjrbD+brb0tl521N4bsVEcvRQ2jUJxtdpZd3CDVuvF
LZFE43tOjiNIazW78w7Ca9q9gNx6rzLuVhLW+KeeR6xcgLaSXI1D40jzkJVf2alY
ru6yIntUmj2SnqN5JvxGDJxJ2J16uBOAEb6AgLI66esIL7sqGp6kdtjz+ETGbH2a
+7A6Rt8SqW/lyvEJ+5TUzwVaWCbdrrFnC89jaakroX6u+foo/PLII+aq4d5IXmZ5
tByUuQ/wr1trj8K4LutHhup+g0eFhMcE44R0c9urz58b2Qk0Og06jJ4qAjcRTefL
jGyl39ecqNXBMHK0mVGTTUwUgAWxPRkYTGQ28Qdbds/ejnvR7/5sJbTCNVyUDnum
0urDuz2ZXf/Df9MnOqYZnKnRVDnQ2YydjBFI97m3jnaxsril2PJsaflTXgxR2GZx
U6GdXyYYYNSi2ieCH/lSYrl0n++9uwDuxH/JazgPzcuaR4dlIXEiakMcEaWYLnKK
WYaOslKP3+u/GxnDgz0n3bxQ+NyYIbuuEEpL3k9s9KqaaSmhZnO6zPNfrwsRYn6E
tg6LBZB1BgdHZi5L3D08Kc0tziy0uemci/k+/MYgJ016UeifM28kUyzCFdeC4X81
Lyzz/dLmRDY3z8v9rrknB3g3V0WcenhvAEICgCxqkjCzyBt8sAgtsyzrvB2P5Oc5
zZHePRBTka5tbtJ3XDQsz8xN6/0I6SxFzpunqhBQme+t98G5EsdHOGeLrJR/fyAG
BeklxToy6f4e+/E79AYxlSg9AuV3B9REux/k9J17Qkuo6XJ9Xl2M3uIwseEXq8Cg
q+Wiube9AktuaNYDAnpyuGMRSxYoSyt0x3d384QKCRvuNvqLBopVW/rZkkSSOLTQ
m+SDlVvCR8lnDgJr5HL4LgfJ5hA9F1E17/KWnsLlrKM3Vp0WcpSFFXaIEzoH86VC
/wClIxybKsqFtbUVIAuKbt+7OLaWRTfDgVgT/JLuBK0KuRVdbS5TUCsVNcLCfNHS
RFy9GWej/cGsxQeXzWAWZynbO/hapeaXOjl4j9LHmdZJ57aXdEDhlW6zLOq+1318
EIryu624rOVTc0t/6muzazarqk576hJ4TiRxVvOeY3+hoMmukvINJFQMCQIAZg0Z
kP5LEauIn9kQFL8h9EYa3QTiwuO4qmyS+Qp7Eycrot/E0gJ3JZOV6vEZwNz6kdiH
xSuCZ2MGuyPDVvueE/OcsyrE3Yz0W1QOUaBNJkvwZJmtQu6xHU1S7XQ6AF3Lii+N
6mwtzaK75QDp3ytMIo7WOeTED4CxwVOvFSAnsgnxJCK6gaXJb+Br+RkQrLdeqCUK
QPR0a1boo2wMXud3fkxGRz2mKo58IxcOWLWlVgbVbvwO1VschDvI8ub3ikm6RrQ7
z2ArQ/UO6fqclJIg9YiBo+l2wIsI97vEmrLV+XtguJjagPiZuuNhWIUesrPdocxK
xUyVW6Ocnn4my0Ag6kJcbtRvS5Ly9koFYv4cPit2+KrJaQerPB3OQYbGaKY5WVtr
6wkAJo49olzKzU22ybprvutuMpC1vn+57oi7hmVQE1XalpHDqTgDY8dyMYGi51Yy
QNy0uWpE778/PjJYRF37ZpRfPJmDOJvf1WHj4yrD5PkPjZjgzyA604V3l2ON6cxO
NAsF1lMwNPuqBAYMajaf4CgdC45fkyAIgYt1R26QQ7fJtbcfFDfBOlohh5I+Ucyd
rsL8OXAEvYyOl8aOzreqOMHNvKmNBGg6cSWOd9CnaCyT9puPURfL+6cTl5k1p2TF
rqG4da2tXRDuJTx3A1bayefGCf1x6Bd4QgyzKtnFd/rPVF6FcCtZFxj346k115AN
kTm23b9sG7ixbebVC67F5Gl+Rp6WyVa5bhRA4N24u8JmBUD9FKSa9D9g+szfGVFy
rTExTZ2yROouo86Ov6MIcCSxQu5iBiVHOYX+Uz0PE27ts9F4/bjho0GLstlTPCVA
zYqeOVzynIjBBHWfozWXck3ioNU+s69CVQrrR6by4ARwvRyCDSKEQraXxgPjo6Hc
XVZi0CgPHxnfaODgNydpV0My0hnE5pxsFJWQmaoNyr+HDZWdg7ia/w2sJuYQWOl8
Jop4Qh0T+fRp+4wTwVBYWG3vbfipGAlpVcUoO1sYsov+liwx+/9nk7LVjIGe198u
bxl0dbqAZAhfqsAH4Yr9xkyJWaC512Zz1DHoQYi1g1ZtXrL60Q0aFNNr4j7bpV5+
PRrW0XtKK/WVN61kgUf5NzbA3Zi7ifhTuXDFWh0apHHkh0PNffYIeVLhCD/BjM0d
s1grQrE6GZo/e2D39VcSnlSi0JPywHTKQJgmS614VFfHB/J7p4pmhprlnWNyK7Wo
maULrTEPZXztUQT91u5AtMRqi+TWF0bdZW2Hk2bt8m4DnOpv7qveSrSB8hg4qtkO
zdJQhBYrlR4CceKkRXjAW4UGlp/AMKjosqCDmNUN0V4q51pw/X+eSgdKq2hS9WZ9
GppNwOPVeoN/L+rzXuXKiG0Q+B0pia4As57bW3ZvRtgo+k3SwK16E0C+J6y85oE+
Qyx63DSPI40x2IPUFVi0c/w0mvw8l0gCy6GBcM06msrBEMtobBedpnZhX72HuEnE
xI+4+TauMrnmjwl8wkOWWny1N2hhBg9Y2dDsGcJsLjlTGpocUXMapNrswLtUmfFG
LaW3hk3ui2Ou461G5dsXrXfyx1OaFiGU9aQLq6CxJkHSeub/kgVMTQO6PNfoHulw
BrZbYFpajEj5kIdHtmntOmmBEokMoaxJn7Kl7InlRu1v3MiwjyD0Wl5KwvOJD/sb
xr3bTZabuhfNKVTwcxFz7VNUW8qcNzAQMBMRSTC5AQMPHsUJFr47RvSj5YZCqxYM
yGgTDNEAWoYw8XSmt1fz047Jho352+2jaD0/yCrX6LIHOwalKMGYN8DM3PYRcfmX
4uZ07aD9BxpbP4AbC4JN2WjveddB8PTq6PmT/Lgbmi5h5ZHQLfwVyrB0vfkNLV9U
6gIK5WbzvmLFN9qRiQB5JfyySO0aVr93l43WWpVX2rF08qJDjxynJVC6nSBixm48
fSnU68QxpGj3j57Dm4Se2wTrechIvpE9jyRHx6/U1uUJ7sMoRGvx3j9b/HJ5dh+p
AxQ0ZlZqYGJYUJyDR4Dj9NWIs/lY+7//8S4FFKNilTVRxg9b91XV4CPlBZVvvMqW
B/dbumx6MEtunY0xgg12mJbZgFwam29W4NWdOzZrwa5gZoz3WFwqF00uM9pt/hsv
siZRF/Kg6Rkc4LsSUz2FSmEwO2cgQxQlWYpCCZYKacn4hm2am45oQaXhvkMhrTCZ
Qn75it2BlYuD5S4BJw35mSO/QcPUS5sLtPKj2pGA6U3Uz91ENS2QDqy6BPjiU/ov
SJJNtdFqM2gyZIMBEth4rVwbbFopesPS71NgYV2063RI/f4VpnKxnQ15cbqOWQoh
n5u4fk6x6asF8YXRuNyhQ7PCV/XnqfeH5BAhn8sMGpHa+luEuN1qePcacnki30EU
8MPFx5TRP4uUuUxqbzbMAv18Wpgrf6xWwAjjlQSKVPFukoxkv5ac07ire6+QksoK
rCw+R6hNmSjVknbSqxBFwlHa/ACwm6wbMjQ5GQporzznXdL7kbdTvqcjmIWMc8PA
Q8DovGDzS+6i2GU01A3sRDuG9Myg7exMiEg29mHuJv/Z+jQNCdwN4/Ytp7LVgcQm
wilkYNq74Z04HWZf377sl+Dfo+h7mZU7ba64hPec6XhJOR0p7UFMNDt21AC6orsQ
nDRuydcSrwWo5GOtEuFyPRrDwhi+CYAaiWDp7BVTwAgrJVEa7ltV3qIW8qowYaY+
i4f886aANeeGI+W/CNiohVxtHyz3JyOLiiK513uklA5Bm5NWImDuz/ARvkpFGrhg
t+R8skhLNluV/Gdcgqh7Zw9xu40aVjnG/bag0ic038PAGjyJxkr0jF1ytxfpl0o1
el9q1GzeTetWQHdOQrnmos7naKkfroGosPtk0kIWEy8QBYypZO34EO6KbgwTQpuY
nq2fL/ro9ojA5krmEX74nTEhuMFI0A0bGH8BrKnn/Li3qxKJ5s60eTHXBJ4CGFZ9
MJmot24zSnUJk2QAtHJ6sTjpLEmS+ZHtuKaAO0uJVHJIZBiCzsqskxOpYFW3pP1v
44vMQ75dRnFwrBv5EjPaaqhKRQDed8kim1G5ngV1EfwW1B8EP2be8p7ieWm0VemZ
j71N6TG7U6s2amlVMPyo/33NjWvNJPFD9SPFQ8VmmrJQWIPZGJ7FclLJBZuOyKQJ
U6Wy/GwTBTRJywaNvlU3v/eqCDo+8DriSwl4mmZAmqSG3E7V14T3yHsqBaAyHcfH
TH2kJkZiMCZw/5MkSoIZAg==
`pragma protect end_protected
