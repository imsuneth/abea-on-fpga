// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:38 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sFfoFhpwHcd9PKXyXMjmH+RvjoLcqgS4zA77t8WqHUNF2AWRjjLCfjGuIvzMPVoz
3e7IUsfWi3VEaumWkmguZ2L/oVuQn6jA1/7PLUj9zvhA1ZLVAJkmexxY4DXvMDLA
K+BPR8WGEWZU2Xfv1FkYmQNrPk7Jgo+k0GdUhDpv2rU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
Gvh6rZL8cV0gnVn6ML7K1wANdscP5l3J9HlBgXFWuUft98eRgp7xp2Zg+xJyXhan
B9wrCeJM/fdpHB+zt+KAivERyp5xTIIGjM+E4tYyIJKDCy/0xnQQT2WFDepga8rR
HFCNUnjwpm72nUJA9hF8Ku1zPsEeGMGdqOFV2tHN4yPk3jNhSsKPmDymW1StOIOA
b5tK+j9V2Zo8Ju8v2i4pWDVWFgk8H4+xBEwX3xSsvNFxRSEg9fvVyipWPVvKffMO
3UiBhnSp1Ki3TAPv9JADvvm/i0Ax3M+HEE8LkwHDbGo/saljL608wK49heMAx9XR
wSbLoFSq1rIcCE4I6pCwomZKe8qA1alZaGmeHRVT54azHxyz5RNkCcYYU4j6ebBS
8nvNT5inGhq8UWP6a51eMoltT7pE4bdS+vK9EXxX7vu+7apRYqcDUJ1T6jB7CoZ4
B8DcVwooBAHOUjE8RdrOT9KDgqZsy4MRPfzUv4eGJqoD/IWBpnj8+wvSMM9JQ6wR
zX4TRqCLTUAotqUQcNTnDSJA2KIjHkHdtDlD2WwFJZNXvrIi+WKCBp2jnHtP5AbC
YpdI3bMEf/4yQqlKFtEJOSVnYIroOGfivOWiNcjQR8n8IesUL36+tdeT6Kyp9NEj
12pqfzu5PQ5Md4jA3ntZiXOjtrJ0wynuSDFubVEembAgg/Mplme0jgElJdM0cqCO
RWKR/KJIN4K0sKxr9isciZ0wKlgaXmzZN7YvO+xqrwtP7ctf5o/BaBqmKIvjtyF5
A6Ip8Gf3JswOXeUpcUm6Yey2CQORi3bbvyQdCDlqQS+rtY/mZencuUs4vhIgyoEA
dHwBv7llOYCKOiL1j68m7myu+/7qzrQRySp1c7DqtUIwmIg9FguUXJnbPJeUMOkE
FJ0kIEffulkvrQNQuSSXxBjRdZfzk9MbwPry0gQIu6CcPrOwvvCprmf+BUf1e32G
FSB3T+AtZnngekYOR3/hJ2j1W836jgG2SI+ivZs2PCjuZVsbS8RXdw+gMTqc7NrP
wqXhqtJcv+0cnDL5+068q47f6iHAE6GKMJZoFp9D3YcLvOLMq7iHXF6HNaYTQATX
pkL3UjocCt+dW9rOx79kbTe9oH6o9LGm4A+Y+5NcTc1oRuWHDQmljoQXO/7nBpi3
Bzd0pKIk8/Qsz9qqTW89aJxmLa2qaQN0ndwkB+6NrKO/+wYAXAFDYrOY1Um3C/nK
GaTi9MAKBSH4+0sGFYQauLxxxzMhNkWA+6nbEa4YvFVgjdM2wllIEcqKWaCKQFpq
PwPCEWck8HczsoSd+fmAhYaD5+qWwk9L1QoH75iVYfJKXlxPaOnOtXSho1Hb9GWY
DTBnPX3y5+AxuVUtsCOcK0f6gG1PzuPpbr9p8uL5q8DfywjrgTq7N6C6/KjtlsCt
Mxz+ljVrlQECqqtPzosXLwNoxAoTO2nkUdPXe9tlbT2e57PEzcr50zWyWVdaaeqP
dZ9+m76r+QSNQuNIy+5k2EsS0XFt9nrpSQPvsVztrldFqU+PJRlwE4pxBwpXFPTu
KrqAEcOAQxeNpP+QMZ+jM42eS3fhJadYiVBn3S+rpo2iIii2zxQlCVuoNwAcM7Mv
HVuA84q7htMpIX/F1Ri/Rd22GqnYosTvG1sGQ2kHdlYIond1OpWR99alCNiLufSM
9HlRB8CaHn1pl7SBq9/Dsza7q00mqKp8HY5vUWYR6jqIrPDUl7l6PJWnjb4GzlXX
+jsy5hJKTUnd/txOZEltD+oidXWE0s9YVFx3qLU/IVG6E2fjYnRJMSmMXWoiZjRd
ZdbSvqrsF/2hD3LmqMjI2HrznS12mIqgvD4Kqw5m/zyxK3cXCpBGW0qR7eyXyi2u
Ihgst2JutmU+6M4YNBNP5WECwGC6ONR+xxr6hwpKTb7mIVqBcFGVPxP4He15rASd
SHmx9j/byHKUbJqjEosL4wqjEbF48l+60IUtu0mBma/BSGI/48/V3prH288f37qM
icRkyEGVBQBJDq//Z54XulX0VpyJDxa+NaMUJF9HJqJHlDAVFVbl57EpQYozgwPg
e2gD6DlnirupeAY5fLvGXjxY0YFa05CdUXWY4eLdSHPQ2NahMGgJa/aoIwTtmVYS
MS7fEojsL7q6kb4UHqO9A38OncBh02JWA4lYBtozTCVCGU7gDqcp7O6Y6NVYZiN3
MA0rS+EruFwywa9SGkiEWSAWw7m2vj9Xa9GOqBhpqDvntPEx3AT2WbpFTD92fY5F
Sd3hGIb4SS5C8rMQHIpDLIX1YnD/I7t2xoNdEWtxx/N5PIG2y3LUP+H3RNgP7Am4
8hhw2WLbST7yh3z0P2HQkXVtNEDIVsRB7wev+/k4hV4aG6zVg6PcrbBqipKwkfMj
mSlEeh7RU+eleA1ZGVnkd+NltSka6bmW3NCoQSgF+V3ttvxHTC0S8QFSvySs4y3h
+rX/bIme8W0ek5LZRwIPxuHzyUo78CFwHKG4jqCgIhydGtIsWJuwMC4WfUhUsgc+
xTnINyUY5t5Pvj1EUptSyi9AQUHe5cEYdoXKWYBXL3uwDQqd+dbq5edrXzEjdCDX
ZaueACJuvoz0tGtd7Dq/9XjMtq+kvkjl3LpiflDvyxj89XA7sSnXzuIdnmS/o8wi
cin2Pdoxx+brK0yhtsAIt+Jthy7w8/BwS37NkmeiueCXYLQjDM/X09JfCDfRfnQ1
zH9t2WF065D85OhZgFLWrVxkA9suHjesPDqnVFGz7wF2ENLzlvgFuiNcoomXrCVH
6/gURCNHyWspQXbWqZDz1dgrwgapbGlayUb+eNtwi10Httl9M9Azby3y/ozj+EC/
rZUh8AieAO0Qa6C9R2fD85KQp5rVUwlzBk04d4qD6XwvxJvy1NOJT1Q4vJE5WfXu
mOZzuC4ypa4luhEO1Dp7cJuUEMQ49xPikbetoHvXjcNHUb62VMoKgRwcgbxK/CyA
OFBB1nEO80X4BNsUU6HHuuK3jWxC9fWT0hIioDJit9pEd0On+e26XMzkbSPp8ExB
79SAmUqw9Ytklz+uI8ZvoteUzTqr67SznRefJnfkbvrt5wCg7NLfrzpZMGShYmqG
DwYcSDik2BlDMWeyErqh548e5e2ygCzAdakaQ4L1K2f4nWC/SfGFnc+/8tHj2V+z
NeuAXsQpZHkOzEbIC8bUhUPoD+Na/0xesSg8OtPH7sJAY66DvjPjGIN1Lkud92lM
txz0vcLkjgNJKXpI/uIyB6gt1md+Q+DJf9HPPzs7iwfzQpoPHV8IyBpWrbfV9S1H
KPKwo4Pt2hrDTzVH8LJUFDXOfJRNlAvz2Gq76xJI9f+Cn0MTzgyI6dgYykc6kfvr
7+OoJkOpBmCey+Yt91pTQfPIZAs7m67f/SZYbbeQSTOsT8rD3OU2QEdTuCobbZES
ATw1VvZ1zJPS2MnGUCSfEl2jN2rV8nZtCY2RgWNjMd7DI9ChtySTlh/LSPsrbkwJ
ncZHltfDyDeLWHT/hlzKEyOtKgaLwugAkLU8wPoQntqj3qa0L99VIjz/busipHHi
uWnBFbr5Ev7gfkY8+koYXEEwKWiO974Xx/3nVo2A4U2K09HcfyMfyPV1fHW19ksm
vkAzJHZr7bvxbAjXxh7LigkgDCuhq8Esn7nd2/9DvqKairA26hrmJsRFmOS+NO0r
6+3xARh6fA8xtO1PtDcclYaJS302fpJHNNEWeYaXfqZChm48JYFoguyKMtsUBrEh
n2EKLPh7qbeL2YxISDsvBse1zRiNwAFiNfLedYlOZKshUOvEW94rJ0/Rypcwcj1B
3YPDdCfgFqaJAUQsZ+MsTDR0MODikmZJzc6ZDDNJ60POn871e8YkIe1JJXB5M5Vf
qdhZfE77rTkgIAMoPiX4GkSpvaoDdIm3YOT3AN9ejNupSy6iBw565pZh4KUiObI3
/Ytj5Ses2q9hkX26+ykM3IqJBeJ2H7C77f/ZGu4l7xWYnMtw1Oz5fBQSaZArrHb2
+Yh3MPZ1Io5oC22LkR1yXy7QQsZyHnPXRfTQkFfgIvIUa2X6H4uhTVAEBWhOayxw
EbhsTuS8dL/E3pZK71t9AvgVG5YFIPw7GAOtY9kCNJXbvFnv8LhLPMQ/X5IEWjGh
rFLGL9T47wxSiGyTPXLfVYVA9cSU5COa7VABCSS7PhfEzzIZMESFB2GjdK535hHy
cTdPfAKnRBJeP7aoFPWhlAPjTMYTznDETreAQ59K9Xs+G+ApkuEKi74rwRGfe28w
4WbCJmV8oR+4oYLnYHRP/5NMEj0onaetbo3lOIZcVwLgCriRAX2d630Nia18I6xd
z0J1Y1IN3+mBmDI+aV8kDtIfkKDMTYgpgFW3XUnRFESrbSonXMissUBF0KHWwO+g
`pragma protect end_protected
