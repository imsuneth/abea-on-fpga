// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:54 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JyWt3AaFmR/mrX9NR7Y8/tdf47aoRNrEOlXV9IGLyPx8pNNx7BS9gF95tvs34uZL
wU6T99MwB9kIjH0rr2BfA09HoG5ELJGRB6EPzLB2xcApxbZIjj3oPD2/FGT62wZc
4ikM4u8q44UCtOV8v+bdsVKKgzEa8C4HHMB0bN3Bmso=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5280)
OJ356/6/t0P6YnjR3c0seFvhdyR2Jk9S5U+maeOrJ3gFlchiPO2cAre9LgTAEbze
5CpPmI6g28TmQBOx29YOxFCyKHUUtQP463bTReofvYp4lrHub799GYL0pB0P3SkL
TweyOILkhZzScYvILDJILtPStU+0YRYEh6rE+s4yphR8IkPgpe0suWPG3fi/dvHc
TJfdXqBRK29k698HL2s8rcG9eVenfJP/omNlyvNy1uYS/AMgF9jZ+ZyJp2EYTU69
GEMYCpn2lvRzu+6+KAL6RBfVpNcJ08VGkog7gwfulwGY1hnfefL+8jx8lJRQlh9N
7ZAtkeadmOGjN9qhMU3sRiYm8BFHpvbm8vEWwkHsShqbO7bctw2wqiw/wZVnCdjv
yPucvGIAnevh306Hqs/Qm4MauS2jXe1i8ueMgFqb5oOeE43AkzgJXR9np9j8tv47
Wc4K8ELD2DGOrlCLew2VGm4xgAl+p2EwXGTpK/jRaj8N+BAInBGlHHROa0UPw27F
oOhvYC5Z9YZjZCCAxRoVQU+9/5qbB0jc0IuXUSLR+z6Cc1yPPa1IP86J07186h8E
oMrok/1uqiGABBXPhRGi2Jzr98tiJ54v23INqVVeLgEe1jdqO6jizmjjKHg8E+d/
XRknuhkPvvaRsRnMT7ukZWpCdlYOYSkTGWDqEGkAKrsDOhl03HbYzMiM59ZZOEpB
/mxGWEF2tgQN40E7YuNNDbeg2/3751xH3g5VNqYmebmgLY8snO9zllik3ZdT8o/o
5luVldwGa/s5jOW4wFdF4goi1RNlJNgqfALvIOy0/aNMb5lQ+PE1UWy1xx2uYuRM
ZCmw37fw2Z7soAGqImY3X2uvGfo1B/0k7Q81mo7E+M/THSvBB87XUlKMD0V5eduF
En6mOkASO9WnqC60ZjgiZ58PL5fIjcH/RcA6maLf3+neuiLlw69Oic95KbEflrJr
f/a78xB5NiWybR2Rw5me4o2njJG1KK2JJux4eidwI+5DBLP5M0hWWrw2+vX0dZaH
j56Ny/Ibt71duyHfQVDDVafc/wcxGV/M8Odih7e8DZ8IUBk/eVC2x8ARYLKVV/Xl
eFbP49JkQx6yjMyOBoCfP7dPI2VNLLN0PAogwiaaZFBxCSrzeB21P/3v4Dmx5o3Q
3tf5F2dDq8zd0NBcsLRJKhw1z2xATN0kkeWS9BvsmeTzDgiQhTM4QRtAluBHFxyO
DJ1huW4WU3Lbz5ji8gG7fr74he21KhLSs5SHOgotI7S1ZQYVYyT3ZEO0fU07xKGx
jWVVY8K6Jk1J8lZ9c9hZPQ6EREDKrMX4UpQumkz3Lj95obMQc2IYc+YJx1q0OT6f
L3XDBkPvTOeJoIPWkScG/JTYcq4t+oyQW3G5C4cOBQbSC4tkXRXh1RBW8YnHYTFe
pRIAZGxuHqIcoXZPgZRcxGlAml4yc6BFiojWmYGwAEafB9ZNA5Z7MVgkxNvwXHL3
I5CG9+aTOjZS1CWIPnBRbWTM+2OQcChs5AWzs6ECFGk4kbwIIOrMN5MZ28+yrJ20
7e7rBXs5ioEKVBxe7xKrN4tRoLuuKbabDXh0RfrH56DFFHA+Q46LfvskHhFxdKGs
VcI4r52E/dpOmJSAXkhiWO+/aDf0VcK6maYSkm2rEJr2J92W2dQH5GquoXdbBXHY
GeYF0lk7JwJyaIFh4+Qn+RbC/u9iDBAkxe3WsSH8cmo6aaMx4oa/Ku0kLcjgpWyY
PVlbbjPF6ddUGXbRW8jl2i2pOUY1etWzZ4CtzLpSd+SrL4GCQksiW9hR/Jv5ZpE0
oT+KVTbSegFqd2vPO4juhN80NL9cNAzARbxD0OG/kJpcUGvi542R34DWLgpNl2SX
fRC92Lift9OokEkTSevSJcJcQQbR6GgxBr10gDwCw8v6qtsCUf6IIcUE1RZakDQT
KqrW2QOOSn++ExB0JRGNCLTz/HPCheYM/XLa+4F37z51Q7ME5Rx3EvHGHZSFUw/u
z4yJR41xGNlMORrXp53G4QQN8mrDZ6iqHhjddn9ZQ/xD5i7xt6B04shmwydQ+Pjf
DYSSl3WqEC63zccVFIWc+zioDT8cVqE6+61R4GCOljEfSu+KgJTnWKO5o8aa1EHA
P1hY1fWAJjHoQc6ZWGcJoLGkzxqdo9N2Lo3xZDmGIiYRWQAitjFkT/9VNIKHdwnw
0Wghe5kTuWZvxTpVcCG8Mx/SkCQ1f5DuotjqTuc7Ck5rVBygSzyLvVC5pSEwwcD0
E+k1cjyC2k2Y3DU2tIxmtPMf8j4bqjjXC9YR3Iuq/uqMNVc3i8tXvFOINKqXGUlH
6LciiYQKcVHreNSF3+eRAOAoiG7NKIuYWx1H7B//KhG2sqBA02j3zJSne1XsN6SJ
pod7k/hOXJuERpS36YaJkkE/0hOo4MzJCSJSxt6fIexNfP4tyq5HqBV2K3Y93yvT
veogp05G8F9UMjby9rWbRVfaikoL7DVognaXRP+ZYpgiBJll0IHO1MSO8KXIsSFG
RnBhQH5Qu/wof8I0vBaSLmwFP5oaSB1wmiwkD9vAZmMdTV7q8JB+GImdtfPJtk3I
cOwyRl+TKZIQx7lTkdih+NrBnbLR0EG/H22Ci1zbsfsGSFhxfvSO7V1NEBWTED5s
Bk/KCECxbvico7zfsmXWqFStVKQbOk8Jyb+IRLSFiJ8xoU+h/zzEHVyWOthS3Lze
niBZM+Vadf4HJHADNArzpjszVDeuOLbyTC+GEZxqa/Bqqi1BjmSrGucA8wKV9lZk
VzvGkpIWEl+kZHswCQhxhQ+j4rDaoo2DM6wZ307hXMto5ovaw5JtQcAPlVpvegvO
T5BsZQ7bbAVecxzCM6AxUe2DDH78Kn6l37XIucIboUZWFSwTROIl+1yN7+DNN3zE
35LHxP4W0N3e6xU6zI7z+JWuofeXWOiKULK0WPboOvWE9JobvuF4EzZX0VvjMcTf
7UaEeu8ozJwb5VoVKdzD1UumGsL4atoPsAyKErMwsTM2gQ0nqyosA/0EKrtO9Ktu
0FKXRNMqG8nxt/DzgzdXQqzQ+l75iJzTcMq1l0h3+eLINara36liujM+37n2c/ZO
kdNW8RCrq6/Z2R5S3bb7GYHace1zPjm+9ZZwvOP4xQIEwvqCb2sJeIr/XQLYmCvO
Jr/BfodSOnrIlCYI+kFg+AVhgqr/Iq7xsnhxolJ0ZYDMEYlQCpruikNl9bforuoP
nLLMfTxAXagKC/ZbDhmOPJuX1McL47VbNxgLKYDcguzF4dDOelE5uVv786lyLvLi
oPYzYMUELEqO2ao81uXy6tlfgluXwQYu2Gm/V6/CCicGEPySJCCBMuFpluANnD2w
9jg2LcyQKAY8sAvaD4MwoZbH2AlqTi86uojO7XNl7MzatpopOfs4MdvzBRnZUXqk
Kld6T0dgT1KphcMMHRznjfPOzz9qTbp3tjFZYDWdTGgJ2ZuYiB2/lozqYP++vHba
iX4bPpyqPQaEhQBXm2xDWCq7BivkhGOtr26cFn4352YiB0aXrw2sxkcNciVbtqoI
KsXxKKSGSodXzrKAOAzaADWFEfuTqkiXj7kzv1YtCtZGAdfXlqwC0vyXne06I5TV
xlobABZB3qzBkj0K8mOi42Kd4MChuKcsOeDM64WAY8fFtoTrmAiZVppVnuw+0ApQ
GnRNVjZFjpectrjAeL1P5zsykja/vRqaqMXwm/U+2WYb4wN1WFEkHg01n07UiREl
hMomTT9HtjVH8prNGGQmbqTvvIMZ2hLaNqcQAijOIFW85yXRM1v0jbeyHZHxTV7i
pAHlx+9s1iRiZDbBIrAJEX+0Q7+xvf+YeaTEoMioZV1KaRN5qnPZRj0WqdBMAL6f
6lYUFBvV1HK7UdFI+Nczper1BnxxAJRhNBwJ5xw8d8f1kF5umlaLkjTbCOx3yWij
kXzEu58ppeW7waS0tnZwe4oufBrhCfHP+426557Iy5hl8S1sLPOJcVgOk9pmY51B
2JpeU2Z3R7zML9iwhnj+n6laWIRbRS2N5Tvdlv9i/NwiUZ8aD3s8QKzEUSrSNvoa
tIAW8qhT9AyCkpTu4gRGHSn0Y4du5w01zYAFigeRXBRc82tMwnQfJGQTVETlxu6/
aw4zs6F54GOYPeLya0eCPH9Q/bnXgM6tADNr72raDPlDNB/xdc9Uo8PzxK1ghm0J
FsD5ePSPtEYGA3HcvmISeHFFkZUnXJSgmBeUkk/a8KREYn0J6HMqAN/I6Z+5IG59
CyJhhPhCHVyM1cP5GIr8OqVTr53+BelNKdldCrWbHQrr31gHi4tz/cKaTlZNPXWx
lACVXz3PK/mpcTXnF6/cXjZ+HcJDrVLXqilkPFVAOH4w+hPiw7RIlxhD+2M9qkj+
ldYBfFpCM5E1IP1W4QefXKnKgbc36ZolNgDsy+UgDsTlLfU6I4RSQdOWcyD420Eo
Lqua2mFB7K87/ePc4gts7VB0+m+1FNoV6YMPA50PaTy3XPlmoHbChEH+LeciZ0AO
pYW5KPTDvci+cYlWtW3o9vJ2Q1gFkjidqfVY9TKhBIvae4NVGSyIS105WOosg89S
YQrSZu9PLWTM5UJfpL6KQK2S7zlGq6rsLfEal0Rd8FF1yyFF1hvboE5FTDJrEAxJ
0WELJiCE8DEOEurYSIgY1PpDZN+/nd91P+ifC20ZRcibiqK9pJeG2ZhBOgRZODYY
QPqOkEYi9phxazkjAh+m1pjxKHkWjzg1rKPhkMHzJtSqwT8jIAFrvKEzm8sDDnpw
onJZcGY2xcxD6nqTsnaBEtMDlDbt1ogc9d6j/r5PpuBlQcGH9Xjyn2jCifBXzPQq
k1B1AkKgnWrqCUAOK+F8B8RH6aGMEaLfNKoCvPHrfYtRUN1rNEEkMh1zn4moIn45
5G5NPGySXg5aml3KKjXEOehLdpmMVbpXt0Vq0fqlSHwusP8erqPG+FjQInTSMn+W
rw0e9X5NraJiVTlsO3arCUvXj1Uo4Afe7FEVb7PLH82eXf9Mfbip6qYhRDdeOzXG
IAvyNhxIjKD64oSVAHZcyjZTWCzjS5bi6EY0zj9PnAwPNsGKhm7EuYcCLxwGJF7C
nOqbKkdLYgeyThWgivVjCdQSj45cT5R67/zYL+eNfrU1hSQFTP6qYSWT1aiwwEyE
OMeTAFvBkssVlnsIFOC0dW0dJgnpg5+w3CYLcX2NdgGbz3ra1zZvGAj28VsLHyfu
8haLkfjD3+zEASZQ2UDaRnOVdEDb9MnHMFnt8FTkVranxSOH3fJoBZGo3cwAAcI8
CeYXTGC0hcthKjLfXTitonZuLtSuagKiEm2M8FG5V9edA4CSdHT+3GsX/vWH1mNU
CTIK72VmViDUbZfAiYnCSgaP5jjgc8EmkanqgfLaUHCbIJRgiWsYo/voyuuNmLcI
csYnjBNMQFrXIj5kV9rdqedc+i2saM6gl7VAXAtOccWUE/oW3Jg3ZgMOXI1Mz0hR
ix/otCwPMV+nRTQM13G3xPcqqtPgGarKkBsBKVa8pkJz0R8c8xEcufCLRyBr21ly
WUY/Jt1WKWBgUnGVNOkQecwufDCxYvszjWHiR9/8KDOTbBfsS9L0IUjg7iGtbGvj
+fYPiXIfSl+Mn10K4oVSCW1zCzkXGbMEfnqwAxHtL71REWsaU//6ZTu6w+yf44hJ
YexthkfcZjOqFaCLs79TT1rmzzi1IfACFx7Aqfr1ObQCzgS12uf8f31Hxna/gV4q
4Ysh/J3zRYfJNJn9x7mFG06NCxhjYPKYahjVFnCLsfxvL8GFqkHudrPMekmfOyp+
qt8DTmj9fEhFPr7phsjxrQ9EpuQM2ld8QwOnKwkm7r24YDTkPhKo30RVsZIEo1dl
f9+XEcud3LojYKwbq8NwQQVkWSa+eykUKj5te2w7Zgx0dUlX5GnUetqZXAoGhEQl
zJ1mCjU+m/OA5oQ0ykYXB8PQ0a9cWL/Zs9IKNmbu2QSlYgB2lymW1Wbbfj+Oi+6D
2jLMTDVj4tfOivPaYgHj59ko4RpT8C5/IqUaixOIVcvZj+NnTNRSpxM3S7AMJ88D
ST6j/k4BsKb/gpr1Tcr4uRQXA6Ecfwh5Gn2SSuIXhdiKI7UwqtFaJ+buLG9BtGsT
RIf34NGiEUhgu0/CW1ZftPLGOJBlWQtoopkKdOOsbdzVZ6oC1bP7FLBFvsF55AEC
3XbIA/cGGbpj+dFsinhCr7+fhu24SeZBxbvM+/JmhBqAe3duqXfNOQYBwLv8qWis
ogyRuvq9RzpSgSGVRHz23xXnn8NfWub3+HkTFJ8SaiTnToXzMG0AUN9z+RFebIdX
5VAGSXA8yxENLF/SVBpxOwqPUa9Y8Z64fRXnvrcZUil0mjdbvcdXhrLoRZc/Zsnv
0WUE+4YISJhEhRjBKJFhaqKDatwUEfL+ExRIklLKBFC7WbLQ32EVTkuwnVvMSTBv
cOaffm/0LmzdM4OQYkx+mXhyX5qyinKQ5QTYO5YUawztV9biHw+3wpYA2pSaJLpN
q02UmU5YFXo2XkienjmvvSVf9YSE2gID/8vfoDJjGD5eR7oRUvEKW8QW+pLpx3wR
j52bQws7DbowW314QSnejEEQYGGLzrtFW7H6awgk4YQHLxOCfOrz/dD89jMi3u63
PuR7OS2r7PQJpyxnE77RxdPGKCqpPlw8a4vvmgasBWI41LSljBL+KgcvGokCgXFN
5+4vvyKa1nH9UgIpvTXm3jOgEV/WuTa6QucJP7vkAIMgwUo4MpOOg+aVsXKpx75c
jUjHAqryysgc2IaE6mG3R3pN/ORpZZm+ZtqVGixs5r4ykDfJNsOM7KfF0dgQu81C
Uk5o4u9ZzQRVe8ggX2+x/Z2HIUf8P5YICFOkmBJMsaUk0DmDXbI4WqtMUY6VxeLI
BDbYmNcDicMLtsFukQXWrmKmouYhWAIIcYdMngHP++Mvo2fuleJ+vsQ6QUDLeEnB
AozkZ5eRizegieqRVz3rExrGlSo5advirvQLcjhKH7OYzGSMJ5mjRVGteYkny+fC
2HJaWcGWgU6f6ArI20Zsmr1SvH+NNUHxMG7CgCcF2nZt9hdZDEdKiYy9LpfDRCGy
`pragma protect end_protected
