// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:46 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PeRopRY0Z2IO0PL6Y/6JvpjUyYk84JU6k8ZUbC9D0WQ4XgZvS/nNqWMUJAsIrl4d
3t/Im9y0ZSMS7KCv93ifbXYsnlDabKKiOKUFEEzW0hqDA/LxQecUosMQtdUk4jUM
CGy7A95/WoWUPA16tGXHaKVTJYcOpi4M8rkZtRPnejM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5104)
ydLua+rWtREOecROiuyae6e25MDzEuGDos3ooTdUQwgGOS9VqPIHij3fDEHG6Zu6
88iq2rYiZhBTjZbLhhmBcFGDUVksrZdoVWtS3vM+6OBIbPdRNkuAbKYAKub7PVbU
+R3gfTLAqxqzHFXGU5T7VmhXGkxsPw2in1QZNe8xSvDextRZ/USO2Grcw1olUbPA
Fg7Ur2nAASHu7xUFqFCQhNPlA0g9kYinK4fcJzfEHR5XKfpszJIcsGP6v0HEpW6z
cugnXhSmkjp9PF/EhLeN8XSxCtYtVmXLFFCFS0BR3D2arP2+jaBlwqFFDFs1i9Wu
MeRphp9oWdfV0iztQs7MhRlv5/ZSpdn5YeRzBZOckWJuSF4D6izp2nPJWzHOOFDy
VudlbMyDSgLWRWCwR1iiF/hvsxLctnJpxF5cScsKMaHF9kl5fdr/8ZjKs7iM01P5
eBj8zlDoIEL8EmpVRdzinMWMtKixArbTD+ar/c2uiPYgpEvAvMOogEl3OccIVAye
d3A0XOU8CTHmw+tkUl7Flhdw1LtB5n5CLMhdfOwTHfCIks3sqz//xWvvgVBH6V3m
PWLQkUAjxDoK8YrPdh7LWbUvIxJmkmH8IPGEAgIaxO3jFLSpzE43gqP4G9uuxrA4
nSZybADPufsAMD+Fh1jbvt5sQrMWpIE/2i3Kvlw5ObpoyM+TQezsvnsjou1t9V9V
QAp/laVIxb/K9kuYp0x1B+LMEUm4ehSsldgnN5ss/N54dmdczQXTSKPlv20qS263
xJFBuG9LecMxJC1Pq4fIrmI4+zNXk8V2Hs9sAMrmEI/9Sb72eUHVLPEftvrlFiBq
GHzulSGu+WyIHE/3dYoisIXcTXp/h5J76A0BjRoEEW0yCU/nmZz6DyMbcCKEg9PM
pD3/idD2LaSHYZCVvadyln+m1/SzYY7X0PLm4XigyCF6SLscMZyDJSn5NPLPw3Hz
ewchdwFck5Zlp4LYAMaPxyhL5GYdGw13v6aBnejHhinoNt7CJvnO0duxJc+0iQca
2z6iw8GDuylbflDImLBVORYpKYqTW+8mp0Gv8UyX9u4q1GUuKhFSNtSY5fHKNmSS
MsxHckTW+gnj0BcIgxzFS66u8uT9uxL35IYUD4Wb0tpkEyak1wPAisWjYnyEoH+w
ASqvon27tlsGkMcvoTewftWMzioqR9T8S7BCm2dUAk6kBLgTkcPA52Qj6RDFURgB
lWCJ9dgfkgQ2705Xk46vsu2UnLbpneEdXxBy4pTnioXBpFkeP6EuMDm5AZBfqngu
3BuXayb4Y6jpBDvLAegyRhPIrzbHYW14585LBwyp2ddgWuDK1mikrpXby+ykfvHf
BBQrVBUk2RQuNhVu6o90Lz8LskK4OdC+4cWBOlHc0DvjfMtWzTBBUaQlJjk0F98h
5Ptet2/2L+rPUqoOqS6EZCZCmzEbn4w5ymWv1ObZVsojal0rZaXjBB5XEzh78cge
wtQz5jJS60MK3IK1B0EAttF+/iZGRBEhspdspPFjBcATTQrXrHKhhefZ39nym7MZ
cAOZLleDLE2arO9wT4m3KmqXzeXsF6bD3TX/KgZ45ik9ceixgup/kucI6B+VevKk
jFEl6Fcceg6kspsvy6iRfvQQ9HtT+oTOp4LrPhWzXB6cSRGcbZJt3BMLPvTMrG2t
fZ0AAeoNXqdoAIQLKJvhJ6nI3Nf94jeOjZRSK6yEFE/dRR8JtAUao8PEOWYzC0j3
mGNOdBLFALOnvrjU/XkbT64gf8tmSSSpJlSs4hjQiHaCriwniD43iP4+KV1vmvUS
USXer005GRcQYkJd8jAl/Fyd1wM7zzY2oZ54YJv7DUCRFAtiJ/CnwlEyddkqPFeS
z+Q/5XdwkDZRGNFA+AOhLCKl4dMAiZqFTSxVRDd7xNbmmsVTVhErydjG0oXR6lFs
RdcEK11hPqlp7m3+9DdHtg94bNUWBBnt6Ms0G3Yj8Ft08ewFw1RCaVYUQ19KOAKw
FcFgMmuNe/zu9vU19dxXqP6Pz1vtOJ/kSgNmH1R2ieQK3g38cBaXp+V1olFbUAxM
0wPvnaSgU5msklCs4KZMcO2QoP9SVZwldLhn7VmGe6gcYkev6HLzpDSEfqe3XQE6
ElH1vofhbTrvrpQnSixSojVmfzdNZB5XoDxI8+TTv5p9TF5/AQ5MWtqgkLTvLele
6RRM/GtXZsbEQG6jCkkna76i2+2jy9kBjwlq70gqfA3R2Wn824J0ImF7p1/ao2sP
JTwd0c3omRkFaR5uLsx4a2v24JqLIXlQh5MyRlIB0pYsKHF1wBm4Nh9Kwo7eANZW
mhGdDUXiMA5wnGrtdka6af/1hLiQfdC77xl+PpDLDmKUjE0qkMD3+zUPmxAi9qbV
FWgurmZNTFQ8OAV7ZXJKQCC8900KnoI9DVXijj8YzRPxgKvEDxmUM/3JMmqK3Koh
L4PtRuC64YFxFDI5lFfvf82iQ7WceIxzp5iWZYH+SmBTy/py8Peh6BID/sKGY1+9
OEbe4Vzeb3H1b5bCBTnIpmUbqHObH2srOLph21ScuI5LVUqdZyNIkhmQsCvxZBjO
X0A7r6VlK38p9LJkvLy2Z6yx0vbA25b9TEhQAzDL9t281hesYc5GDuj52PL+nGp5
Gm+pb9q8pwDTXKAReUCOFskxdIBLl9hf6d1udKML5C7wGF56EzcsWKTpi5cFDIvN
YpvyaI1PsGgLIZ/qB0l3mQrRi2ocqnjQpwp4L9qcrDo4OTHLWZ76kCbQ2bHxEOjg
JwhuV0JvjJ9uFKKbmVLY8N4XwBmfdoUsV1pR+45n5S1l6hTmlIZAwyE/SsEXwFOi
UTREyUUtUy2gAxL0bT7SiQ4MiQKJgUKka7gut721C4QH3xGdhisuARXg7nc2K1Mb
oi6Krr8z5M8TBg78UKIHTfkCb7tTBGtCF5WH2GKppmnMsVfiQkLcMyrSLJDAZqV7
je/NMir5FprxpCiahTm09tt7WiDbTT/tp5+15L4/FMm3I2s1HtCnQkybOpX8jg3u
V+pAsvOp8MtjVU3iM/SiNcVnPOUk+08OPfJYDEfKQOTcUYigLTF58IkqdGDDjHnt
XuTqaUEsIz2cWu2FynzoURyMNgsuxbpl1DBwD2RvzqCoXq829cxvU8ZZvuIRDuAq
2FCzV7vx0282LTD3fGsiwfPpqUA/psECQlaTEdagmIaZpaLocGbAumKjefjxIieM
Qu4K4sT+qZ0j/F1u4rdANG1Dua1iuM2mAu+R5HzhVMc+IJaI8u1+HjbT6BGkDifX
puAqV2QjaODA1VwgJdlYjHqYUxgdrxt0aW1D8IrT2V0lIyjrzFf2IpENKHeCV3Uw
t/plTi+wR2ojpkbITu9Z1O0w6oDLuf5a8PHmuq4OSpoa+Xj8ZjxlsZ6tmAzKliaM
QhYBC2CpKvDc8PvMY6F//sBa13fggjpsWj9jG+xN4eT6LoEyhPUDpWLaA9S5sqzU
KqzMquRehBM5dkKwXe4HwbDt4NWKJVp1GlCEKgr/4ciBdz/1krsBEoLMOUVuxagu
RcebGQYLGSHRmr2rVq8Kr1oo9RC0VIr7V3cJUMRZ5O/4tItmZoLbtk2Ob9OLyXkx
iITx0InBtowwh6M+WSSJoyI5sO2Xi2h4i161+cMuiiUBcQktzjPQPhGXkV6Qfx3Q
26HP0H2N8zN+TPEg+qq8m763J6pB6YFfTRljS8VvsyxmUl8sO9vfBfFXZ1ct/rVm
OaMjut0BdNMpwj4rQobyrQS/5sTQGLUjDWRDYBxAgbwa1nSO3ifH2AE9qYRwdT40
PkQp71ou7ORd9zwH4VLprs0WCz20vFUdvUnaOesp9mp6fBp3GlEinKUsB6pyceFM
duQBDGz73mMtWwCNhtFfjV+XhfT/6VjMYME8bduxX7w8ehXTnyxgY3YX6nb/Kst0
5vTyVT2OCx8yEtpeKxnAaLUWUP2lLUdqfNSdkaGcHON25ieaief50zHqLhBqN45a
xKZZ7YEAp3kABVfZKZkzu2FMv0O93YegZpKo4Em9gt2vSP4s5tcXp+V9k3TyUT3w
My6rxcWQU6xDbJivOyKC5AonYOizYDLr3WPfjCXQFBNeJzTxDy0ljCa/9nBt+9yx
IHOOIg5WAcAsYXQibqlyDUKrQ1GpAHCb0AJR6J2GPQJnb8EKgjMeRECmiQ+00dlp
CD3zcAIUUmXGuF9Y4uSqiN6N4TJqOBrZBEuH7h1cFo4wxpf/2PGsyEPkuY8dcq8U
y30JGreWqCaWMP6HR6/g5Ixhr1JY6VcPbg+aE11YMTK2Cu4kTVQInNGnbfG7vCNb
mM1ia3whL2T4avVwFppvxa9IVtjrYm8d4n1NX6IEk4ZmyJJxzFuNyUClzHlBpmvu
WmiGxKhbjcawfEPN8HWteqC0pMmrqP9nIt9fPDQMevBNzPEfpzv2Ufmru6k5aqhS
YSYC732Pppfhvgb6zUNeiCnXEEVuNFsy2vJUQZjE+lv/eCNji+MUCDFf7f8Zv63t
Ew98D3LxBUS5wCgzYh3f1yE1kbX2kSfZqaFXjzMRYSYZPM1Q4n/BR9YUe9Rv03yA
uCdH4fh3mb3YkVmcnq2M59vPsPorRr52xj7sckoyoOnJjGBqOgrJEAqT+AV7ds88
obh4Vs/85Ndu69iN4tm+t3aX1z61X34kg95Xg562YY1tYqkVag66ecSTuoYbl1LB
FcOiAOAbOETnVpYLofEzZLV233Mr4jizhhSHDdmUKdSeIu0nMWx55fwxFioTzCuS
zsqyKguRXbbKzcJvsVduW7W48lFKtwsb1jluJlgwwhLLP+jkQs6l5M0bUuuohg+B
2qh+sweC/xexF2ehi0HUL+TWON5fMvgkakq4WUCOZ13P/d5ez++5AqkPCn7hTP2a
rui9vcMEBJ2g5Vg5YzZcG9lkpJ4DaKycaSruMbSdMKDyYFWYI80AyYDJL+SFIY03
XpiNNrm+zxhijU9gr45uYu1TRP8PWN1KYVB7k2xdV/2nn9eZ8mo6eMtbGCYHPdro
7+HoQFOwRBKbaQHH8ZVCQ6S/u6IOBnaERlqX6LF948oPL6Xch1pxZM7rpELchBQ9
IsW8ZUZ1t2Dc0UwbYPGipA0PEs35cw4nW0kNmXQr2WzT+fhpBmnzGbc7ivCPqWHZ
Vm/jhU/rV5dQC9RHkwH/dMJ1EEfKq2s4MnRRcoLxONwDTP/EFECX2/cONzdUulFR
VLj+pNZnpdFcdu00rLFqLyQxThjpkwYrQwxbaErLc6/r1Ar1UjLTtHGB8NzDOE9d
IVdXP/BwqeT7BDIwN8QvKevzmNE6XgoY0NRdYkWDH1eT2hWUWm8FYRjRpyVYkOEH
RpUKzfXNiHviXaEhQCb248t1He012DjeIx1JzHR0k2IC2UTdot3MXmqWhSfTRzh5
q3BFZdwIUvgOMH1cSgX7vyUIGQPPQO9vHpQsgtFbFEoItRIg6bQ4g+dPN+2iURuX
5Xq9IsNH0L9zHQ0w60PU7LSAwzAEYLt6NOefQCBvHDmtiXEdjJl6BogRMJf2+SlM
YskAZ63WxvJ2VdKtBMOSmkmUL8teGNStM7D6dEPqMS7FbPR/von4DCeZ7YQm68/a
iG6NGcw78x4mMFy4+XSB3DXZve6XUvzhr5MIAu+sF6vvlbfcan6vJURdeC4A2OPG
mShNomKzQjFVb2UkITbAS2MRrIlDTairUH20osqALa/M6nznJ9NiPx+QazfABi+M
cfu2xwTRl4SrySsO3Jc76yGDR+Yj34Np19PRPJBnSEKvYccQtQVrfC/1b/V4NlPv
yEqqS6cvpto3WI7+DWQ3X/WI1xtS6oy5G/TqCGaDWNIiV0Kw10Cu6zCG+uEP67AU
5c0FbYFlvrjTmaSgO1VJeKM3kHBoq97Rgj4ZUuvZB16fTgIiQ7madx5sABHJRt0j
eFNsIbOaPj9GUj/MLIzFIeMdBtNA1miyoTfkQOQ/lTC3JhSJ7MJtEooTyXEfCq+k
5dy/u4LNXENhI7aQKo38eTQV0B7RC6brk4ogL8zY8asifaUywt33it7EdhOYgu07
ENC9OANkw6q1ua+G3DseLTIqTXVX1lFJa8mQ0qEDpIpbQmbM++6ZXYVXmXuilq6H
UlrPqOK39M19bX/3MI3T48edOvLorf2XxylZZ4ZnYfVITblNKGmyEnbdvifgnmat
iZMLD+nLcru/1jGfgYwePW+nM5LAQ9reBjdkEer1u53E5DX73KIHP7v23vMj4V+x
hpiuuC7hGERc4ZKX7OUP8uyjf0CevSv4digSlOI+wxiE3S9DVweF82k0CMpIBN+D
U66IC4D0V2io+t6j2l/8cAx74Drh7v0MugMTJg2XPZZO9Qr4fwSJC1I7ho+Yg3IV
pk88tx6oTM/wP+rgGtsZGjvz0jJBmszed2n19hQ6Wb473g09ZugfG8P7FidgJdN7
KnYWtyZuz+wnebanx5c3WOGnK2EVWJXE4QcFw4lERpH1sWD8k0yJxcUax0mzlM8S
QrY07DiSj7NmBI3kpzneQovi6ekGt27bPa7qdwWmewJPdP8GnUe276XVk6cgBk69
9dvDWa6P7mLqJzkfcu4uCH4J1hHoIz+8j9yxcPoZMztoLvnWj4F8Bmztvk/2CIkx
dTUDbCEAPVMWRECABRvWi0zj+rBzN0zvXtj0CYdvcguJJaLDdSr6RkCGNqxfcVL2
dZuiLbAiPbkbx7gaGkZm0y1V7qQQ2C0OJTNq9ZFomNe6PYklWd0KkkFiMrG6jQsV
OgeJrTR8qyf8XXMn95giV6t2tiFsb9KF1HPT79GzksZfGsAc5Hv5L2r7Vx7xJiXs
wntwY1gcERunfNbM+/08rg==
`pragma protect end_protected
