// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:55 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MWWgqK1K6rNKMFI8Tz1g55MXVfooprA9aPeNH63WJWJa92YQnicNWvQgZqqRfrwQ
2phFOgPNU6sFp1WHe0LZDubUhMQeUqs3v0CNC/vj5IzwcPbd9Woj+NOhn8bivjMy
VDSQVb24vZYdoeYzxP3u2T2kxGHmQtKAuvS2HYcfO+Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28608)
QMSfjuH463CcdAcztVC/KZQdv7JVqSqIuJb9jTD4xHZM2/Ujn8y6wIP6bpmUdrhJ
F9PlBjbdoYrBVG1nyzXsP1ftVDS/ZZMVVXTGZQDcpxJXUvfdWyZZYkPwhv0WLZNM
LJ+tWENRIS/nytDDRn/fjSFMzf4s/XqzqbAO5yTBCWj5S//Y1bpKaZjpedWAyw+4
LYHj5NyZyl9o5df7mKo3NScHpxZ/DE/lfpegwKz/SkcG7KDANpfnQJGwk/Mm9RDl
h+d4yyQoUSnwn4IwhdXrSk8WuGH0gHngR0+FSZyvPOEUpSmLCHsTYXd87ryEhp2n
sqMp3prX0s5OZhzjfuPKw7MAf5Pq7r0WCEWX+lIUMZBGqkTcXW14476TkuGcUJcA
Wy9sC2sZ6Clrk5QAs6lu2G6oqDMCqVpDqD1gyQHonh9lVBwvynxAmtrIH3BCXJpN
IGbbgcb0jUYIzbMakehgY8QN43A1Lnf0i7OpIDHHzdtfRd4ztUc9xr6C2ThJwy4J
C2zbQpoMXAL2d/xFvEaxgGOZ4LZkoDl0cu/eLpIsmDHeoibPYcMsUYckb2zaZe4F
ERCkLfkYRQFSlYQ8JVAeqotHedJi6+g1KaAWYOiooLJ4ELOOeyZKD4Z7R+mB3U9y
pJYrAaTuNQvXIKbxFjqBx14Qt1LjZhCvNhupsEfMGfYxECtaUAsvBUTEtprlJKK7
umWfZisI4tHslcdftCqIJKHcA6SxGr/voiY5H70mDBFz+9UqcZWr9cGEw80JPv5q
6IzwcmMoy0u2f6ejOIp9v4RUGaK3R6AU2fqLO7EjymInjfck5s0aQEHjgLMhkXBH
3HYpneHdA1QgMgcMp8IXNFPtwtUWvp1OhyT1oA+bROsqf6aKYYrN5llf7woY/rWk
idMCh8K62Iq+9jdRcfjWBe9MFarWAD+hHUqg6BtxiweyLG28yJUMEL+s0CQYwfWk
dgLH2/iuMfobQiF8NPHuN7q14TXyBhj9BFyathYUOjEFmRtALzkplOFZLxojdESc
XRak1OW7NfFLw3ikBfd/FiBp63CSmUGPHqARlaVpLm109Ls7VzUJ6ziVO3xUoPxR
YyxSMfNNA/J8C38a4qcATKVzmAecB1nyk5puYdH2Xn3yzchvJvbE5lisT/KJfI6E
ReCQ/pLutyje+qIhdT1w5Eyu/UgdFfaDUrUXDvz1l31YobkZ/navhNtIZwtvuMM0
MIgJuzdnaEhsiQCLH7zf3XLI6P3mSy+Rv7X1dqK8pFh6U9QKY46nEzd44+i1A3VV
kB2HJhkwcb/MN1CW3P95IDG1hBKJMwicW7AV9qVBj0Tcu2ITHs+vHDFx3qSjy2I+
W56iBvwRL0ZLDENjIYGZQPOUkgkaBcX4DflHEgAtSTwg1xJQS21euxE3x7Svg1HH
yE4oO94IcTUNWb+ovLrKddCNGAXstg9JhluUP5l6e9oWas307vu3OH8c5NU+1Ifw
yQSbULGv20AMByffHIybNQmoEFSMhMHV2cPan47wejUIiqYt+MoneSpFoWc93CyA
2/8LWwp0ahk5DUx1LKWE099M0R1buDuMC3tJ7ri4wS3ONynrNA+hnxOJR3/NNbwk
9gmKDIts82I+CY2ZFK50iV9StZFg0nzpyyykzaP7PrWZ+v/7KfI5kKqxd2CokXPE
EDH60bGsOWgUvb9+4NNFrptDAOBubFZRlhevwDDf/zP4/xJ1dB1Vz4K+WZLSy6++
ECM2cTDknFhF8ALBua30A4hsyS3cMmuHHh4uYTBO02lCu9Rdtzzg9c5HYn8LJM6K
B0nnjaTdRkAJrfVCzBYOIbt/otGX4Y0eREQnHtRG68N2IRPKmuNOAg9mNLLp7ev2
6x+quied85nHwwcPHcGkpESAjmj/FERVGnaJvBu/gtwEEcIET8KuzjSNbFHQjc8O
P4tJxGDUN1aSfzu8m2fWW7xjdxeJeqw2ZMm4YMlIY1bk+L0FbNeb/JF2hKXGd9+f
YzlUbzcUN8D+hbiVGpngNHXRcoGTDRkHaUL2wRPjMK7+R/YzM/Hz1aC4sK5uxDGR
EwbXeikI+0Yx+dBaLfC01nw17+D2BFocTCagE0FRnmKyyMopHjj6GMEDhfgErZSV
7L1/C3i3Qbndgw97IqwCcyynkWHEzTyA8H/Ip30mOcG/R81IWeF9BZ1MXY3ezOQs
LKEqYypxYFwRVuqn57nRO46C3WQ/xt6bB+41NMXPkC3XV6YliKtK+t2HqaYetJ0P
RGBE7ADbE0XWqXDn/4ja1GxX24LZLIsLpoO1OzIE3TaNnETwmPzdYDEsJGwv3XsB
dGeDUwAvJKhhYs3DhCzAMuYgcFBa+Edu5mD+Rff9VzsDtq1F4ghmqybEXR/V2RnH
O3dNvX3OBrq+x1CGnkF+pH2Et3wsGGVaKPVve0NdiMJzgYZ82NBHf5XWVBoyp/rP
yLiN/azuiOn9FGzkLcNJPshIUAjtMv8rW9FNLserOH6b97UmFOO53LvTQMF5Xgmy
lsMwi4vICwpq2mSqjouaLve6GDOfl0iZ3m+IyUi2lREpzQuasaHK7InXbmYEUrGB
FokMIeW9xnG6m2ziY13Su4kUwuDl0Wu1f9Znvihb6XlwpWQlkzqcAYM2iMFtgG+E
94up9YLI4OOt7SzvVq7TqqvlBG1fZZHrKsUVfGeTqZkZeLQrc3yoNBnNow568DQe
F4OIs7oEwEbC0lIMdtpuNmexDbyvRlCltnOOW9m8Hzocpn/w9w9gsQMnaA+PDAMx
wjNN6SXoDkVrU70HfNOheIMHPAix2uqZrJK1OgaXqQyBx6jIx3FYmDjSAWkxNOJW
ITeDqWyYzOXeznv3iSg1/466mXM6dNHcoosSHUYlAe3z35n170OPpreZEB3aaURN
Zwyx7xeCK1OZ6GzFEH+Saa/lrJ9zP4Bp41tcPjT0OhdLyMl/wm4ceI4Lh8utTMGM
a2elpZ7y9WMcBKknaUiYxvELTQ8xjxaIeFX02/Cy4pmY/fuz3+vA66zYq+P/LwD9
68K4yt5gE16H0CZTSPq3nwR/RbnOV1hlzZzWCAR+XaTzcSeN3FublWdgbrxNsn/G
x0R+SYwdub+8L5rmyKj5H0Co5tZ4IpxMoy8N8f24BP3TtX6yzLYQsJmOD43joJz8
2uqqIXAA4L9WdqJZ7u4yQIvC3rQIMhHAuy6YgHxDPNY5YQFafkm8F6N50FU9vAhQ
MuMMD94g1RvO8A8krCDi2c63216w7ztnvmGv05Bf1giUxK4byAOdvonJzJ6HVN4u
ZoJMLe9DSaFkS0AYrVFeGwlvw+BQGgNqOHjc5BYh28sqlLwxJ8giMSwv8aGx8NP1
yBeCnlQ+/y+6DvB8CrzBJr9mD9m+lDxaRWQyEHaI46/ZYrPIDBLV+YgO0KjBOZnM
xD6wSPUc1Z5P18RfF1yDt7VujVgxnK7qK6Z+HF3Br5lGYFB9d9VSPm40dYLZIulq
jDTqB+6MembHiwa4tccCGZIHmAodqb2MC75BEjyMaD3ceCCdb+1UbdnoNA1ocnCt
2BqFqbl2coMWhEoS0Z2+zbpw6ApZyNfkQLaerHffQ2ynx6trsNAIQjSryvwx11MS
mIsHI+RokCbO82WloyAwWgGJHsQ/Isv0qf6YdMt2AHngSt2xzmkqI2ocjhWVf4rR
BNOm5u2Wlm8QMRJmqWa6kluaTapuVV7mXSx/F6dagc88j3zxKQThiMaiNyKiUANg
RsSVgmLKZA/sKNji/UCENKnIKo+O+uCPuXnVk8EPgMbd7xWNfQ457U82efDVTqNG
QXWOwneCjkEt5IuTXJtTS5JKDAXNoqna05F8ZQADT9GqZGsaYYFU1sYeaTVqmD9w
6iNQn9FLCDK7y1onoKkj7TRerCUM6vkx+G1gz/FHdq7YlUC/jAG7rrBQBAMWvFZN
9757esg0ZxyBu0DcWoi0EzmXoFl0d/WJWpuc8nfcuSKmeXE71ihlxayndJ77mtFQ
A66q0LhLn0uM7G2M/djgUwd2OxpN9CROJPcNs9EfP0R77O9HTI8r/xGg16c6+uyy
/T/vNBUOCPaA61bxJB6z8vVRqydR3KykdR34d1tEhLnOu8nr8qvB1y5DFRdyBwA3
OeOli1h1GnSidmpEpZcpaCCHmNkaDCi2OiiRKKmni2mNtx6JQb9+KRMzk7yEml0c
YPl5c+BNj1Xfsg6YdM7CnjkI420dD5asw8Rtp18/dl3KpJIDFAFlIKhrXtYKtEzz
IqDsO2HNOL80vdzA1gCyXPgH/ETqwqffy/k09KgdRhLFdKcPCXhCfptGTLnXf7ie
ZYKJxpGjCqE+bBJawev6UAwqS6mdCHRQx2YalJIwpCdK2cECw0HpFvmQm1Edpf/7
Ppe1zFuRuYTFoQtBVNw7AcPP4k360v3/fxC2Cg3cWjvKbLJhB/tj2HwKLhhriw6b
rNnxDLIGu+WZ8tdHJ8hO33u8p9PVpt+jVLQPR5IrDAPhb2vlytdzmUoESu+aLNRx
3ZJ9cChPUM1gffKmPDAUUiFxkQt0/IxG2MZ7fhFVSDh9J2JsBmMmJOKXrAI2tedI
njwQSP97eOFt2388Mj0Kfy2Hj28xhHS7/Jb+yqadLlOEtHQA32eDu1blk4+YhVB5
ka0DE2j3IOmsgoUd89sxoeKUpvvpYFCaF4anGhql09Aet1q2cUdMJtgNt+N6k2/7
JD/9kd2UXQm/cqxA9ZGN2dyqEIZXOayocPS0RlduezZg5bCV64HtCnGhSbS/k0+5
7J0Hudh6QG9LvUP8rleHYMjaZu3PLhmUEtzHCBzTv7YPlHXmp29vc1xNC991Ian2
pJAIIubW9qKdgUzF7E4UZvGl4U3vZJIZ8KSa+CSqTLs307u42rmha5pLGvDa5nhJ
20xiGTExIAJLmTFMGTJwwd27T8GE8sBr+i5Qu2hgROv/NFwz+bxXkPKF9AwDDciz
O/fJxFe+TS2XDjcXcIQeDGcpp/ZkIX4jSLYjgi3a8ATwIHAS+suqVbKfjCS2X1Ku
X+86TZoywcQlviQTrbXOnLz7lXTCaZ7GUwcGj7vnvm3XJNWINYUKQxw69LyI3i9W
7wJF0j+fJ5fso8PwIPq7YaS4ipzLjU6b6i0Cib4BEAt9ZbB6y1lEZ7zrSL3VhgcQ
MZMVv4ossqWiSPk0eI0WbSBOBQ2LOAveDYWfsTCk/TfC9jLoBRtpdlsCmiI21fZ7
Mk8VutbpygbWTg1vRPpvRnSQ2Nj9kThDcHRvzUcnBepLES+eRNbqKl1TH+8muvmo
Mmi4haVttl1oxfYFKG8Ln3rodgR/CFpC45jGjIIZN3MZgoTztVW/QLIKhTErNY80
loja6xAtEv0RQl92ZGppSHnNfXLr7l6Ci7lC6Pw92vkx7pwHQCfCl/dyybub9B/C
jwf7OYgIWZ5eH9N7KFk3pC5lA2bHe3ttJtcdHuvYrscJVu4Z75ee0GKHCiZDLt3l
7hBSi8p9JwXTazzsZZxO5i7v0vJyVpQCCb5pIbGWeGWt0MNz5RYabOTHbqd1gMYZ
nEt1308OX0cCfl6xMri5EDxFhq23xoqhgDnVbpeAmwlQ5ju9g5rgAz5uLhN0Z6Tj
nxblLSEWZY9Sld6aSy9bxJQTdUgxbvHdFKDG3TLnwh9nXF9qIdMIhId9Om8WTtB7
DmdQhjU1VJVO3wR59oauKXuByrXExoDh3zOLUf77dZa1xIfOKR22cbF1cM2WFSaT
J9ZRkB4iJYV8ukRHjl2fg0LSNtXRmoUcQY6lLKhDS8We/e3hoLsW9BnHHjynj++v
1zgmvCMANv+a7xC7ueIq5rU2hviS+zxL/1N3kRbKRRLuaqICDtVQqGlUWF4y6m3J
COVWQvFk7h+tEG/I3rQCXBdsB9vjo8VX9iYW8GShCgnGMi5f7hzoi+sWncBJhTmq
PtohJPZMCZQ6J1eH4hRtoCCxqbOZHNa6T6lRlLlK1XIFt85psXXZRJ/Eeri/hCN5
uoizOhC5DvJbhQ1GLXraIgnUw8CdNYpNOISb/Yum3aqlHLMZaF97g0cbwWWPm2mM
P+SogpCy6S71JEU+2s/B933Vl9N9bA4vSnIylMGIEh8ITshYcUU3Um7JXmCU9/CQ
W7kmm1G4W4WC21eMeNPFowpjauGpYtMxsh2X9H6yizP/1blYs20jQz89KpmrY7X3
HCQ3CXIKrjVhHewVp5fFyarIxfjwnxO0jUsplmKx8b0DYEK1ULH8pIZIuvaTtXAR
xMLT1NgxWJ51dQ226lK/SeHf9nmlH5qkvWOnWMFH7OgEbqB7u1hjn2eSs9onFL7v
YzBtfnzNFWeC5bE9IoEI+c1IW/KM/g//22FF3uI1Rn7YhAfNYMTSA8CA6HhwU4gU
sxbv+XHWMpaa+BHQXat6aWkFrg2FLrZUWoxk7g7oU5VU4KCbVzayxVj+kxE2RD0r
M8y1HTvjfO+CbQNj+X+/t4KV9DQnOcAYPusaTUJLAkj8L3fv/EtHlwOdjdJzyZLs
TmXVVFMZBqjv0msOc4I1mdL2Id21hgucDK32mtnI/HWlUlEN5PPhbAWUNFCgmhwI
qxIZPgfYcquNGe2Q1LajQ3/xYppI7T21d/3g0sCBNnSVT7iL1yk5SDmXpu8Fk/+K
0wPFEqFrHRkkasQXPYg0u3zHyrxm9gb8DDdB5Uf2yhEDC6ysi8RKUPOXmZWL8CJx
0+5ubsypMX1bAQK+zC1TRvGbDAILw/JfpkuV7x8YOpYqFr9Yw6pu9o62EFnRE+Kr
yPlCMb0WGn1Ma6JX8fDzokAihIPk6i7cwvtbDhaTkgU2DwPeIAxUVeTHxurwofbc
SfrKPF6M2bV1PysE7f7NzRCbPXnOQJiTvOu0XvOXYs62ZKyLa2e7/BBBBXkENftT
TwVM+H2Q+sRt+FoetNOKO3PMBCxybdAmLgB8AlHgsDZN3DHybm+UvH7qrEkVP7fR
Q8C7Osfldhe5qREBenl1u80YtTdSU4fHiFXxjY8sn9BQ11Tx1BXOttU0GGY7m1Lv
dquxz5Z3erAWkjyrs9YoQMKRTOhIG9xhe96auGFTA4YHrxG9tf3O5xkDcvPa1Jvv
boSS5CXOZdrQhIdtgkNYyYahmWoRaA7goSeKbpzdig2/LG3FpC6vIvLzWwtVDAR8
bhgS8Fp/jqWx+Lh3p7yMUGOprdYZfeQyHVTq8/dUziREtW73Gel9Sot/qy1/8OAw
mWcEwjfOp0cUz9FJCbLMRcyudVpSEUdVJJYP+iMEhzN6vUbr08EgvMWCNkYOWaBf
7I3KINDU21xf7GqxeJx+QHaVuMHznpKKckclbT6nMChT3A4c7LwqPPjGdcUk/HWx
mvqfrUIKvGAjO/ex41JcSgx5AfsL54LPwmAU6Plf+DWqyRpU+lz5wbtyCh2CQG15
pVefN6ZG1GZ3DJtQIc0VWwKkma22AXHoWY7qClVoPRc4cwn8FOtVL/w2Ah7Ybbf/
Tk3P49vf0bTTsKRw8L32QXZUsOKu2EbmS6CD2lX2/x00wkrpZ0wUkVs0YcpahjOY
DrUjtRXiF42qksMnUUCM+X9ifbku1iIV1B02teGrzwcjxHsq/gqgJqVYaqD19qLE
SUryCOTRNxh4/mdJgt/c8nhbNJbAX7M8bntGFf2YUeyKXNIcWXDq6jrumKchYpq3
wDE1hS3rrC2Bk6TuPzmUuhsEutGd23/ImlKiexu0a9KXvaG5xUWmybufnBQ2zV3d
3lwb4QngOykwc7iskm0knhfZqX5aT8IuL1B9SpoPp1J3rwXxRW6PPCgImO+DXKs+
D6Ot06VCumbQOxTBoPhRot3rbiVZhfTP1GPHq3SzNpF4yWJ+23aCpnpQ59k/afqe
rjyc/1CyxixMYR/Mo4+9C8a1+f1b7xz/j4WWunpl0usJ3jAh5Q5kiQlDOplH+5Xg
9vHpvQvjvf66xvFVr0bRrNWn6vuXC9oKMdGOo4I6Ncjfhcshiachbl5SJo9Cs6sk
8xspVGJtRHnWs8TS/lkRiwE88WCbLtqCH9sMIAijdu3f1x45EBpOpU6KR8dzrCyN
1dTzzxXO49u6CFSGPjCHH2dtFSShNautPh+7qwnSQgWxU1JM1enJRTYQbXBXb1E/
Z/fHlYyV+wfmB50Yxeyr93Gc8PL1UFjgqdRXWoVJea11pEfheRrYhJk33eTtf+XW
ObSa6PqLzZOmyhgh55P6gTwhAmFhFuK8Rk9NC/gs3DWVamHhSrj3E1pILBytsITA
Jur5SCjWP3oItj4tc8fChgEHPVvCmlmCl/N2DDQ9JWKc39XxlLMhZBmol4Soi3eM
kesLCrf5LN8UnoC6q/ISu+HtVllsnPD540IU2afJdZ9I2udRLIhUIR8Rni6LpQJd
XX5OnM/4SpVajIr4GkzU5gKcstNQkhjz49VQ+BLx+wjeX+O0too22ilD/ZdYg+CG
aHDHPOdrkKCeNVPNUr3RnB5Dwlvpb6/D0Op9PloHVetq3PF0T689+dJ4EovpUwAW
ZY8cZSuqXrbVKIbcy94gdycvfTT/7ZW6oNZjW8LkvP/Z8FK0VEKJgB7Qw78aiTZr
/WeFxK3ds5RQhq+2VTD4+E/G3TYl5wM2mv6aJKA1aCB3zWmsVFFsWTNFjI0mYVL7
sKwSRHMSsTsAlyKF3+9ctBFmBMaLvMs6w+GWNyZQ/kRAmAAMMW9OU1HKcZMFxtZR
vY+weoYJcliWECmowDi0MjmxLyzuSRH0gtbYz2UGSJcswZ+3M8TE1EDk4htgMuwy
WfyyQ5qk7gFIfgUXiOoJHDwzZAPa+IqUC5QjNQKtjWcrGgKHeNZSgOMK/xAQi9Va
SicCerbzjZqU4txHba0cQfH+YeyJMOHlFb0TF/ZBNKBObVhHuvpYghQbS/PzjzEe
Uo/xluDCKEulvKdfeB18R24tjShj4dq7h40AimNmZprzslCnXskNMR3RYyZv1Jgn
XKJWa8HapKeFTexmgUEAplYmhPcyQ7QzIHHSZuhxjylGPP0oRNeojnwLCezdBJGH
wqTaljyrBgoklsIaR/3rc0sMxaakuN3aZ3+FvT3/Nd94mrwVF6ffEDdXYYVXrX1H
kXKjARm5RLdDtadeQRWXLFRF6js8vlWKvUQzq+CSWQ5b+AJc4EDhmGCAV+qa9smF
51LyFzsFkdX0awO++sY/fw0S0dlz8cRSyQvwFewqSRDWRVWpflnrxl8fc67QJ3FS
n2Yzbg6lYOhET5K2470t/zyae9iGM3hMFDpovWXyHhdX8eJgUcF8llpz8dkqPkei
I4L4h+ufKfw6HcCNrLTG5fpzgPsjQq30+h3GmOaI0Wi08kuX8iD53Lh8q7F6cn/r
mWKDZ76GXiPAfgIpJbB5yvvx9OtHoUTDxeeOg80jf1y84NR8vD6UbQMcLh4joCAA
EM5KVSKkElshpQb2F+fa5kcxciBYMzQNn5bPP/O8Rzpi3gPkxtMZ3g5EiLP8dLcL
5sDS2rjwjGr2HmFw5pwhZ77PPCuIP2k3JFTXM7PoVDlPxNyKnkdiVHMg34seiJ9c
3SfZZvrrqKCA06VxgziW/Y1Mu4ED5fI2HEZ64gQ3vdj8QOmXoqyNb2CuPMVAjDAl
hdnUbaXSv4iqx1/B/BOSH5j46rD+CqIX7/MrpCqWitsS6XRixmlaIuuUsZxYk3iV
rFH9ph36Fra00MHXZ//LNj7WcOXDliJMojlvjtkZqiYYqZMaqKWeACBaO5Kz+bwQ
hxpqy6cVD7Tk2Sw0ZbjkAtSjfl+epGMsLskLtnWG13K/fA4ECcG0eMlWB6gZpcLI
XL063GQCMMftGv8uT/W/h26CxvXiLArsDNYbAg4CZn3x/IGklATXInq6m2ndmv6c
rKexNdXXg5mOfRtX9S3vd9vNNrrAowH+ngS+cALOJXvyWJqNudbHCoCexIeRcqFf
6/+Cymh/boAsHNhd1HUGFR9g5t/tV/E9gs+CqukEn2Nc7N8Qzf2dC6+PPbcUaG4W
KZvCgwxqNaetMVbFqzhhtuJdMSwwPUkJlw6m037UQs6L+Wb658hmk7uub6Hr8Moz
tyICr8DuW1FOJCNecmr31cGN58F/eCw0EK0r/3n1xBnxq2QUrsmM8R/PpNLzIj4U
bG4CPJC/it7lX/pS4U32V2T54MWzEvRu3hMYllh5mJOFkNbREi3XN8s90gVlSPsI
jAqPTNK5lyhBG3kaDq1AYH3GH/0Ui2qi6vhpR8rZm7qHVPbxFgJNIcy7E+NtbyPt
K/xs3SElIoQE1DweGUzlOLXAQxXvIdmjK9F2zZD8X++YVtpApF5kLCGNma4id5aa
kdSXY37+nQ9e00FqO1sYJ8wmNhDQufYmYJO9oKhFIJAPSGP6OYI85ZoHxKHaDtd8
y5GrzDLSYKLuP0o+ePda8A1YB0nCGlGKhYdtBtnk/PcKD3QQNv2DgvcU/foiwZeu
OFz5Kujb8ka5JTSdklr8nJKFL6IGBMqFcjCWNJRdDF9BjtdbbqoyUMw85v2/LpE3
62u0ickyVoo9lH/GD5bypLIOjj/R73AMnjaQbInuS5R8X9MOOEDX1MPdb/4vnlqF
cnptWwlHd7pXDxr730upgtmiLamY+r3FkwnlrksI3U2iSUcMANgBByiKOfM2zNOb
apjJX835CCZiTYta9oEa1nWZUiFxbJ4npftqO+D+qUQ6LJ86Uv622qMy9mRGsXs4
osCQZJnDXsrWo+Bwtc7k+byE92Pt1xnVY/QaeKUcS9nZiXDoLG6T6a2TYpxGEWeS
SfmQl3l1rzy6DCeXRTxNT7YrFPQOyPB8xsR8QkmuPnfb+GT78sTi3vhtB4A1orV9
aakfFsrV+NtFy9RW0VrF6LfaWaxIuFjTSBiDKQrHzuuCqAhtaM4zj5rOBpIhNltU
IUku8xjMg72RYzW8qVMmFOzvP/R/5UWSUSvk/NxYCNR0wsVqUz4cuZSQJ8LLpQq4
fP9IigVFeTQcaspxNorwNuNwyty65FAl1P6Oi9kDhag444dPxVbQzT8F+ztNoWB+
o7lYEVgMfv6XEmCsdCcdSAeeGYSxyxA/xGlK4bKAikNlUCWeRMbbRCWy2zRR5XXr
XOtdALA2DScnqSP8uZwKsDsY57AQugY6rnSa6IKWzLjAOHWmLB8sAWsVZ3nKGz3/
DFE55mI1lIE1tqZdgFV+yE69oV6gpeSt+mBQ01gESrvZUMLcPH7mG0+LkrAlIPrI
Ef3eQu/OpZUt/MY3U+PR0GMpiMfkUU4JeB0mDzTFbtStwKkMDYq5nnHPJpBm6GIa
e2Y1zvPBfHHXXYytngcgvCaW2Wt5iEtzM8J52eKxZU/4FrJIndPHn77ygGEdTNmR
ZUNAmbKko8Q6M2Lpz9/xN9qmyfmHI62S4QHSciFcdFobcYXG6aika+r7qqpsG1Hi
3KiVkLKpdZFOUj2JEPfDLK2t+CcTHNsFk/ez50GnLhw1nYnf5X6rCQexgvj9ts8J
dSRAWWgbckTpH322WtUgueHFUt4Gvk54yRFRN3xX9JdB7ef3Xgjg7Xbpzl/p3uXC
OMmYRXnYecCGE6b1htbBzXgUTDi17FFn7MLjI27kUHw0w/J95wa9WqXtC7ljF8mU
ENJE/gx9vJPSMK+ULVfeSro5YighK0hYcLKrLBJWT6nYI5qHSfURHVZ1AoH1I8vU
rlS5a5NdHTsWtiuaRL5nY9PFtheWsQGwqHzhBL5EusWCkUWw//8Ms2SiG6ilYgao
uCdtQ4zetKT/c7mlZFTknJjgEC41TDN0rZzSBgwTUcb9MnSo0rZn3pzbG26V/qZX
4T7WoN2fes+Kkni8r78K7Ks2GaQSuStPKmSlqlce9gvVgEvHWYyOCTcqpHwnvpYK
NBPiMamvzYiE9zmORMs58dlG9IioFgfmFJo+U0tWCV1vSabRsre6GJjgYTj2h3Lf
TkoJ+MXGWGuydWpOmvXeA83ZS9mruPnP/eXJJE9oCizLOxHQEf5CQYVXgnDxwEi7
e/eT+gG1ujMSAhDyxdOAz95VX1/HkIip3JPVh9/zlHrC1LocUt2kDSCOwNlh4jJp
s4HAT4AAGG+OtIVSZLnaYnttWGE6ejg/VIIy6uVV9r9oKNyz58K19jpaHjLAKBtJ
ecpYc5K4/rPs6fYmBLQYWpb39vJUkw5hmu7i7EfiDRF9Qu1r4uXj9pS8Z1RuK0Rz
ZJ3wWuLp4RxBxQxANRVFV4Hx6ddG2R3NighL3Nrcg7dD8w4ubG3ZHEkhIGCVBdNg
OCm8GM8z52L60CNcpu4+hLCkcwAfPU7VAlhi9uQynL8/VCzRqKC4UgnVPMSQ4UqS
0C2NvzTIZ75LCtC4wdbnyo4fPEjij7VMqy0v/y9rOObFoMQ85Yhx0eafVLFNdgS8
rSfkxOUZVGs6Iv6MMUkGVkNQWVU0SufyX0gIw0rs3pxTk1UAL9aV9biX+cMT0bL8
DU2co555xo0yt4I4RbREl9s7EB19G8FQNF6U5ogLRMxx3ORePV+aE7BcGseubH4z
P66yEzP2touqIIz3NArgGmTmTrKDweKxUWzRf56wITxyaZhsqEUZFT7yFpcGzIKL
4ziX41yXeR0UsBac46UfRXQOaicbWtQ8EJ6qIJEEUXJZTVQygQUZB1/oQzQysW51
CWUHCiGYV40I1YqDqpsaLohES4GwOtq2UlAJTjCumrwteqkAwTC4ZGwGc4a/4JQp
FTHUjj+BzeVQouYNJ1S/vuwM0GN/sTejpRgNzGdy54UWUK7X79/jQkLIKLHp4Vbe
vUB1NyK5fwMQnqjC/0DCa7tCyyiLOp4wUGmu4su2qOnh9KxCrmJfJikvDsCd+1G3
+1Ej2/gvkOFMXsEaubQiuaLsYWkTmsK4jx/wTOC2EhCvr7773RENSr0wC+8lyDS0
QkggqeGD/zad4r+iVp5HZeYuWC6eLxuqpslUKoefMbjJ1k9QPoT9A2X1F2qDrZwN
JVFDwNh8Cik865zHS1SWJ9k3jVv7huW699hh5OSVYcWqGCKPTrjVxmuJ88z8l0Mt
SO0iqKjFpLeXFShADEB5cGnRWD3Ccd8bHA2cNsisB42QquiktW5+t3g7XJ5KjyOC
RaBisFv1Hsp6ZxocjpHc1Ja3mgxHL0sH05bEzzC6e7SAP15jFDdkMwOO2vsrPlCf
pAOBrB2+wuWmQskYvLkR6VBKiU8+NfxCKNzyn5nbSIVOCc0EYl1DWrg9EvphciaU
D2lZ1tDDlkXCudBo9GK08oZyeHkDPJF2ab7x7ABCi6fFQuJ9s8vyCTB6le2gq746
8pVFotbspQPPtqS1n/C/9NIliiNARxord1fgMMgGMlm7YNK3T2DGN7ymkRIt9mTt
XCwI3txRPi4wOt7TM8Gko3WcoKGky1kceXpYX4qNVYSuPCdVPW2r6IMeOjT1xTsm
zWRG83gxjOix0WU1fOf5xHycBj6oOK3CA5TkA/JLBezhnTXPjD6Z4Bh4MRxgF2Yy
EAOrHVoGmJzK6gXzbdAt9YML0lyeQDeP0fk+McbeVYez1czrHB995ptfFSmLAtMr
1Ohd/s8sC1IaI0yrH/sUrHwePaQ87GkdpjGo2M1HtdStglHLH/QxNCc94kYSFCnn
aJ1gcmDG0eY1VvJcZcntp7xKgtYVRDZ6QvO9g4pUk/bCDSgFPrVdCzZxFF6QBib7
7mjIwBqeNZLK54FX/RyJTO2alv1h8XG0EUqtRJYwxDQbMHoa6S6ilNip1AXcT797
07uNH95/DZC9pG0Edo8gYfhiSTa5Uhh+XldG2ljfGkJmHdUUzgg77vDTD3Y9RiAh
RPY0PdwlPdDxyBg7TpOsMXcP9P+QTypRXIvinaIGK4Sok8Aecq1l/iKhWavoNOAl
oMgJXjss2OfNVXQyNRavempLNETY3WPsK1RvGG0gfJ4RJQkWAntHpwPLVmy3nkIa
fNKooSOaZwh+Psi3E6SyZHZWI2Es6kORm2JfY4fsJMczrVDt3wpG0fq3P0/O/Tao
I2GWvKXwya4L0yrofh4mm6xStUOEjhUwtbaDXPZAOqkYXwW61bmCoHikCaFeb0oi
Nwq5p/5Y5rwIYtOEKk2i33ad9rcxEcezSiWucLuv4LIyljqFqvM10ofPJO4ghZ2/
YRaZYcs2XPZU1WP36GKF3BLHaMt+gr3PP2dYAE3wVel1734TjToPdd5D2beWhCnd
QnwiXn7xmq/8/Okj/KnM4FA/NzLliKR/prH1zcpuGBJL2h4/jqwe6Y5hUFvn9JtF
eUohT6O2OZVGJBzy82fPJn8LyTz8SWyvZmRAQz5SZTStFwMKsDIOTRHXPbQBcHkC
VvzOUhxhVXboxDGkchHjMk7VuMy+9CvX0OHuZwHJGPUA25ofAIV0Hl+MM0Bcw56W
GnclbVakAFxZsCTayj3rfXRURSpeFNFW10nsctKsmiTRpw+hFfq6l0KJHf37jcsa
Iv8pmpBSALPwlwwqHfR0cTtl2XmRB5WhbfawK6r1DnGZM+nxgTt0yeqsXt+U2iL1
Wl//lqHpkBiOXtm8F4c5C0mU6N6mna8ubcG/eLmazmBh24CHi4Qjz03gqUQ3l/tV
BUm+455eVX+wdCOcAilwWQFOThZvZWdcTC8U+yBrbY6vegWzkqaGcSDUmN1ECU1T
Um9RJLIuntBV2JvIJeu5DvGFUSESUTauRSdjigkpN4j51X0pOfA10L/CCc34NBv5
kC4D6w+YtU41G+ABIPmu0fwW5cDjcLVuph7o+WeZwLvsfrl+lJpOWpYWHCKq7Z4a
HEoRIdesJ9TFPq9aY/NuucRkCn5b8EYjANfqfD+mxa2JMmw4Q4wVO4AllRmX8qOG
O2nnq444j/c+c8+PS2hvLWLS/n/khhBA4Xk6u3wYPHmhIgvG/hFC3MsT2uZM5Xfw
LUElyyKLns2uL3QxzEkfl8gP/JF5+G62Ou4+VwzmNUEODtsu+IDoCbo6QEL1MVJB
lguwDrKlQbcQUTXL0qxt+lOaL82fi5AeOm3BEJaScsi+28rj1wsnikzzFQi7GL3h
Sws8mgrndQYebaoMo7o4igGjY9P9WMVLwa6o5ZRlmaElnTGI0RYW97+XLg3FkC1e
L4Oki/7YfjvyrcIGlRH52r6LFdUr6ggqAyKuRHP21VGsF1oe9BZXHM8PvCsBfYuN
8nPI8HeeC7RQ0DCE0cSTkvVPSBuwqDr2KYGl7nORGioe72r/Krct2VgNsgcMemUz
83eBV/DnqO0rB70MCUwtCve6z+ivGJr6p0YHy9ds5SmNha1fxZDh/LzoyKyV3PnH
rPHiLrlfGm2CljmcRJ/kxSbKU3RQ4QV9FyotmoRfCLWiEh+Ofz++lEIqmQ8zpWfp
BzIO7xuRwkctHbn/jrFmreHm6rLiDmnyTMjy6j3AsZFrpqUF3qs/IWpUVUAiXMd8
hPrsykLJQBXqMRUN3+kbSnurNlfTFIgr643MjtXgzOaigyn/oCSF7NraOa1hkmSi
txjqdncdH92r/12WB+QMAEkBxBhygmIbhWMj5qVvGeLiHUZJK3BKG9abztbGNEPp
Q4UUm051Dvzj6iE5GpyzeU/zthKpd3ewcY5+bxNh3cRn/atrFFeThoFknEtbdFPY
uB5HaGT07fGmw9/lxlPmGr2J+WwNQ3m0966oJX4Zu/+jDfNhEJ0PzCyYoeL/Td4r
P7/pQlEh3chBBuokvv1RpT5bMPuPHGraTlFqxJw2huDdmUgRp9C+NmL1N6xBr8w7
zCtssbLuJW8a9DwaPNVkugKLmx7kOeggBg+jNdSQwoStbZRr5dVQ63VF8HBcVJFN
v6SlrpD3BifNsCM9YnGIIJ8TP25e+9KedTrOAZyMY1bhrX3XJ0/igYoR4DO+gn+I
D5r7zsnq3ZiYjMZ6p6EVjLp2FNntkD6JGx9hZRxiQShmzhzcWHY/KnEQJRC082hq
VT0OeeFrqgB3NwePGtxkz5lLsUwZL/R8MFS9SGR4kW01lvboqYK03HXWEeWwWkNm
PXCHCQ1L8iy70WQIuorBeHasZoRGYYJdyvonaOooIQUjuia3oRVAXZqdrVKpjQb7
iJNJMOd3zukuR3M0hFlZdr0UhZeZalUdS2OUppv/+gTWaVMpgwy8rEB6RVgpFR7C
UdsocDx8IKjKaN+fbRB85k6a2gTzJgrxl13KgSyh/1OBeN1A5daAa0I/9UhZLbq7
Htr65QDZWK9n918A85+u9OfsbYA7oUuML0pGvGr569Ll48RkxpyDjJxO3lvr0x0b
/Zemm0WRLdGfItOJ1shwt4NW+V9OR5ZFYxWFLS2Z8KrSzukREdstjRNcJCvmUkBY
5Bo8bbrWSzov/35zbK2Y4QtPDdsq8Kn29TYBHoe2QZ0CZ5POBZyiG7tc7qloOEla
txoA+UHdhOF2eDDvjhgbPUdXFX2jU4a8Pk2rs/N7FmpiPWFuuJ65oCvE+Makc7iI
2ek5Tg2U3aiEc2ksmtUpwK8qxmqfVrv6a72wPVdCgLDDrrd6l2/HcsXuv+j+3qLZ
bnTFAPGddZvISZR5yFvlETTGlQ1QSv8EJ5+2zzugo3QZ08Cx2uHRjTRg42mLzxvN
jBhHSoJUwD25d/o5dM/be78xx+aqaMTNSFu36S8idb9Xov1bGkx+dXLXInWz8Ufk
ad5XHP0Rv2NHQruAKWePER/prghIAH5xed9Q0dFMCo1Q0TgYrIzp4fsqiV773nhL
8P1NiNUb1Zh65NwKKb08P83YCbloYCd6TyjhA7KrwFeSyIpswkw1dQarwgLHDKh2
bCNOgb2s39+mejfXaJYj3NZm4DloJ8Vhek2EfR0MDn/hDaa5qXfOhTtg0AfRFeSd
MR1KdXtEZPvJQ7E7f6dijvygawpRRKT2gDpKhOtcjfEp5gj7GI7F36cdlaCSDgk7
LWEi+6ypeYH604qo4FH3cvx4EUKAcZJHJBUlh0OhDaGjePWPeD06Up2Bv0BVJr8E
0knZ+govSyrDJIIHtCngkBedVvi1vsFM/Qg2qP2/OV3VgDTL65yJWvuEe5udYw4W
TXeSSA3QkwzeGYcmCV6WYtO+hdJiCMpNa8q0pCYG83ssVS79+7ZppMHTfV4FZSxk
y5ifhQOCeXMbNzi/OxRciPJ2EZaJI9BYyJL3p8hpLt/+i0YhFpiVGnOpPRB1dNQT
vHjDD7pF7fWnVnauG27dx+69DaQJVs4r+9PfU7BdgYEn8tSO1MQ8mFney4T5S/Us
PLLIRtZ81QzcmpXIT4WJnGUTrAutdm1hWNyJNrxNyN7CLOgLQOrLw3otaiCaw0XG
zLWbr6MsIAUCRlvvjF7oGW245cAL1PrvJz2OMdc36vkeaNjSjf4wjOcpuN6oQCVu
7GUo2nf/91lxQvC+WSDlZvrSRO6CzWw3FdIxYD5K/1QPj2xN1ExX7GVGgnGN1uW2
SUTZP34GC+cdZenupcP9t13x83UCwWT/QMOXrUCc0swfMWcJY1ux1DcCn8NnzSgU
CzFcoDlUrNptY5STbOzTbZh9IYbIWtkq/DYMkit4udgY962oCklTqDz4ui68Rhqz
WQoUgsCJVjXm8stN5jBOy//hvN16xAPrK6pyJoqIMSv3DFn94JIdGvQZVRkOd1eF
kGPb1dAaRuCAyO/NykBuxSrReYYMsL92JoJmT+CXMQ6/1v1SFzPCc0DU55nS04ct
BlPIXlVEl3i5qillgWIL/BEMnq5cu+8/K+vO8poOcE0gdBggvkehA0OqOwD46jy+
EvrVBuuHJXO610ktgQ0hF29ZkkUP6daEnHA+P/MqffHcieGfDo6tO12hERUJee22
m0HbolFeqSEwSDHF6Kgyy8dqQ7wCftuUZfD7cQBbynAjkJnzKBAl0p9RT9BwpH+O
Zk2XEjwDYpPM/Di/r+8rA7pp77bSbXIp1BznFZMyQtEGckE4NkmSd6VHLBA5SnOH
ZgwoGVtO5MZRhjB11aJHpDeXkmldXIDHKQt2ARlW9OiLIhC6UcGxvQUyZrZj8U1t
EU70CUcw2fBXqdOsqrh7ycmfNHA348j68B5PlSPewGN5q7VsMq2peNjEv3yDmCe1
P8cURTdhEO+n9lKaVuHUQIuub1RmZns8BOrlgh6fra5Wrmb5BCm6wYfAbUvdDoIp
NOxes5M6W0dr2u0NCjrkPu5+CygAYgbi6diqIHEvHf07GHH+HP6sGrrVeA1uOmjQ
ZiWK7oZQ0qVWcGci+bwMdobmKk59m2shLG9j8/T3+C67zq9TWVSqSF1F2EJ88Md3
VDxzFu1Kz+nbiZ7ZFZRQJjwA9IOdLOVSy7if8YZyYWAfeeQlfCjWSSSKBFxWKEYD
HIEMSdquKjoyaEPQM4Bikd7Wf0YeXw7SAxKBpzIAljUjhf7N0FDm49xIWIde5S+u
mh5oY3VBUsKOX6BH4EtqyYS2jhM5IiAl2sgjzpbpOOniM5X5gyDFef8lz34ZtNla
cFvLeLocC/ya8uTFFPuwLUnbFThXWjW6oqp2s1Kt8ARHMyoPnaaLy6uysTlC3qt+
+Vm9Rl0W8AL4AFJbP9uJMu0sOYYCKBrXYMSDF/KMiMBrOMti7z8ujphkPNZwrNzk
MpKOUmfaYVmrU3oNiIVQwTum+2Hgm/TKIcMOlqsSnSppG0anY3TJLtUM87LKzKMq
lnJOZOwUaNiyNmX9MPNlDIfUbVwyKJrjXrZhWafOQ3iiKKpafoaikxXABwVEMwb2
Yh4ZiMEXe7H0PNHhqvR0h9LmE3+7zN1LUhSla3BBhCCs3ondiUPpup+qtTx+ZEn5
3WbhTWW0kysYzr6eM2eOIDPpnhdqwaUrCRbNzwDiRXdoaHuHYn40m2c/TexZXyp2
XcfG3nz+0pbey1tz4ES8MRzrYYsd6zFsQXvPC4cetaWECNHprQE+Eq40ukcXL7j4
6Uo9fZHBqLfjUNWG6YTKxgf2Cnu2Q2TRH0odfQfDjO0gfDyhxI6JTGPuOQrJGLOk
EW2kW/twfOrWtvd70O6XMVy2hvGl+faBKnPEmsS+/mKQc2VDEfKMTGPhDF7VtRuO
WJkqYmpBPb36LjK+HaS1DOvIP6byo9axC2DJP81Bjqs7BqnUpUzNOovcOZ5A7jwk
PBhfJNrrf5iEetJDnI2o2nqqjT1rGN0EvJJ8oEA7T7xrgG60mvmTJLi5O2ahQQZY
lGJB3NuWIibNp8guZ3/fz//plUNuDylUgULSmLVWtQg5qjxFjz+XqzTXHfG5PhSF
oT7l/7EeuMHnUO/wXkS8FSApiKKYE0yA5VFjyvkqp2c87pUujVE4KMERdyKcSUhu
4qgLWxo/43xw5uplrJPxTrFau6lStE3T5p9XD5oUjJPVEvrdHor8NnHxcGHhR6Wd
CNlO99ydZgCwa602+R5jw9trllOn9/5kvvWPFdcwSEgVzL102DQHrd6N8fN8OxZs
TKmVOyfaN/nZkXnbG4pBLLe8OEfmMPwISmysXHDlRHrEFlh2LC+vCBPC0N1FYITi
RJyTLXKWWQRk+jV94Qdg5Sq527s4P+sUo8zxUDeOC1WEK6z0qNBPsEZg4WLwerpN
TK4qBB1VNyNjOK8JGtkWsZsKSTmX4IhZcM1ed14aO1y27hECA8Gk+7gcrMm1RLog
drlVRh3HJJtVSBaHlEY9H3tNvT4Mog/vG7M7Ud5UztlwAfHR36V1qWCzRbWsM2MI
LbB6ED00QFZCJNU9f92eW51d2kmmHoRl1Cwz6lwuBPXN6b+9y1+/dRS1eMQKZsYi
RgknnBB+6AklSBzY5TyB1a1qR0fQv+uRNUyiiKvF8we6/LUBMJazGy+RyNkGamcx
tEkr5AIT0HqNeI6BjaGyAEeWJTRQUAfpdgjqBVTOvqN+VnYslnEZk5kOykKWDMc0
FgD5hgMBXmo3+u10UCVXEIi/G/VpvX6zUhW9oCm5t60tkAHmyt/DlQ0Fzpjma8sm
dv11f9zV7gX7gtq5IIxwjQIs5M52gzg2GsAXE+qSPXTRaDusSCudO0gW/v/+bBuo
JoiMLKfioRcB76d4EJAyfOQDMv0+oAXAnHSmcduN0zpxS8FGw+ypvzu3RgWfffHy
QK/p0A1fmwQ9VX9tLkad/TJwAVYZz/CJbqVw4DqIb5n3e3UOzxshdhdhmFwpUuQe
ri5efGU98eeF12IpnCNWc6JY9OLsboNXrnAPX8pdGNzAhcLkKdeplsttKPw9WUEJ
ZDP9Q8ZxolsVMDGycxEIaptH5T+BLHs744nCcLxi6O8oh/L3zFoorQcU3a337MNA
EB+rLCCjeL1C9P8zke4CahsF7zF4sebuxGuAVQIWy0SwY097I3wN0vEYnjg2rhxE
ZOZpL0sTY+585TJ5oPEn38/QpGOzqQJpt1eTVIk5gX0QGqGKcnJrHxxuvUcPliNM
i0BFdluPz8ou3VtXiIWzzczVUhP1Nvr/8Zl4X57ImrNsecjVvvmpsmyTByGQuLJ5
4eCmZjOq4CsgA5K+RHB2OJIjuoYnqxGoim1LeqKisOxGULhmhb8ImYS0IU6NrZDS
BzhuXSiJvyPTs/Op9Zm0Y6uvbVBvvmQWh35ErJWPZJ7m11+0aws/ddS1JE+0NMNG
KIXXeUrHZq45IC979GXCfZ66rLHEgpZ4ldBZxOew5SNEfoVw4OVZNFy5tJURY3jv
APsJ8L84FkF6yJd65Kz3dMAk5Hn656m2IRiMxX1A8PZW9JCx+SH6d7v7psIgNYDW
7wBeJVYd3wVJrq74CBpwXJr5PUSZtmvKqLOVYQPBNr0fDEIw8pLgj9veaau4keo0
3x9XyWzije7gLfs1eknBrgx+w6NNRDSbOs4pC+T49YHu5boHHOQe5dSPkfZEYfzj
2AuNIK9o82kmzikndFBNUtXdVzocmTZWM6xHm9C1I5tf2SyKFsXyWfV0RImQOx+C
ZYTE8A5lSs9kn/8tOKLrbW3Rn08sDOuydTmdeMhChb+tDkTPpaDlPWZm2BQ8eYxn
uWf8eHEPX4YCoxFWn9W5qh4xZJ+Xe75Rlnl7Nf+O+9vXyzxi6Ki8bF6kbrtbkYL4
u/O1Irq9SvyntEUG60dRSUQal1cszRuBHJ5z1Shqxjmit+KkQP1Ec+qM8EMQHRur
efAE8rt/v6GoXpTqdDLI6fvAwbeDVeZkhmbjy6M8s8IbmD3EhsW73bM3frb0Lhsd
zPqda5/wPnJkaz+/jJ6f1P/VLyocWkvTyhUcwH/IFh2LRkUf2FXhXudeTOSrm+RC
aNqDMoSReRrd/Ls2H68ULIbB/+2I6uTHZBLB5yyddxKIita3WiiX7XHCm4tiq3xP
YDZA9SNPA+aTMVT/Yfns+iLDvOCaWSSOvK5NLlHsYl0O9tw1gjwjtNYdPeq1liAE
COfbFe+aeJnliBUjV4dWN8hVb9ncqtARYlm5L8gWEgZE36z7swqKVe+ZWSv/4xLW
66T5fLx/58nU2/1LhD+hPim6sc5FHQs0iEJCZ5hSvTW8ioqeSXYzqP4Cs0m8nPN6
mkgOs6+3wea+S0TjxbINJLo2gFUsVxwhj1U17CdxbsLx+B2aGDGgrqJdM+peYBQm
gSMn4yUNNrE8QrPLuL6ln1lMQzrIya6zgXR8aG921RZnBpNal+0uh6K3hD03Ixzn
5lgtfP2L+HRUaL7ov2s67ydg2w8Mouy1sFFse9fy9MRQZWadNIST3Nl8v/aD/9FG
+RYhgsnTs6TDJcAuTT9LYJSe5ir8kfdx4snhJamu/pDSQ+A4ZuS6HbKaZdk1JJPQ
aLXRuVDVuKOVVQ60rnOCmxsmgsndKMgJPFRMnifIN488luHp25m6Zyc0sj6sWQ+d
4eJcHZHICETHAH+bQTg9aJzOi38GfIKVBCO+3edA/3kuByj2VGKFBDC72pLJmao6
WFLByPhDDE/ay2Rwu/iJI61o1CtDnvA1rwYfIOdeG0Udx3VcnyQtCHIol5pDBz1b
ebQt6LP4hHlizDKD/h4814iqQIjIR1A9+MDLDptINn+nvIffCniZ4qAt7X5FSH30
EqHpcWH/TELFsOe4F7jFWiqBhD+FuNRXOT5xIBiiNwW6UMeWGneabDBol2wnhvdK
qmLgrv3rdWf3RGX/oebsOJOEDh6vBGrYR9YxQxZcVwTmfl4JIP1wSXOW5Hw/+NhO
fAaoQR3gaOWYkIKymckxPzu3/WVD4hPb72AUOPn0ag9CY289QWVkrMu0ycytrOHY
1THG5F4cvraYBXlB+XYD+mHmusI1Jy7t+QSJvsfFCuhfa3G8JNO59qgInTbsAsVL
WWMtqb7DZr2MqKEJbu20xkhGZtU3H8fmBJywDQ9A/NxiOrOCylAV2veTGkOtQBWE
JULEwDmfB8amHcW6QjOaIbgLoS0Zp9bz6+7sVGMBKnFEzZ8IEc9//K1M8tO6pti5
+STQvnPduwIOLeQZMjw25VHWsYapsXpIUnlPik/c3ajuHs6vPgzRbAsK9OLAHjg6
E+/xVHNMklcTcpjgEKwRliNC2Qf/iDfslUBqk9M2EiHBQZfpwjQexd1VT8nXPgvU
MGNjN9x2pUf2kukz0BI0siiuSa6sKnG+m3aC/H19k0MH0WVx7/VAjVO5ieLlukdW
iZIHhGdmhvXLBajB3VKDWIqwgu08oLQVzIc/RxFltmWxtm66Rv9f24jzACOjHrHl
+vkLl5XJHBzSuX55ubPMJI+WTZZLTV9TvDh3SIBtjKk1tvbPHeQsVAK5mqu/6nCa
wKjcPIKnU4q3OCdSkmYe6rFdtVsaI7q20UX2rj9RXZlSgMLHC93/zt0UlBKEKYM+
8P0aUj4M1ZTuJk5xgKg4c4GmiNL6tsnM2tu364oNINcXoD5ywJIwkGVRjhVL27cx
XNgOa/sRUK+2iufreVvn0N6Msz3SKu1w9KHspLP5VJOOTVMAnog4cjmRFfrdNG4+
9aBCv0SDpRbNwc7eO9gzDp74uCF6cQxQNd6JcXrGeXRXMoBkrtKGaDIyzQOumB3t
CuRjCtSpt/AB2fbS1MkcgFcqdcurfpSWGDZhLuLZDUNqtL1oKIEfBuULOO8HOKKo
9EH3CyRSHSC/kScBRZrWqF68O+Y66/R0rn86q4qfF5dtle/9AC8P7rAfLbrDW3ji
RXdWCj0bu0KhkrMThZU4ZZw48UHndquPVAoqjY9qaTfaj49TqkT1fmtV3rPD2i27
eDAyOsuvJNTk3VwF2q1vsfVxMslP4uVrAgAR33AGrOWgsbB/SYLaTOsF7ENq3e9J
/f2J+8IUNgqwVTX4k/gBPGOM2xiHU0JIHfNiN/khvSFLBunVoQRuuXlfOOE4Xynt
Eb/9Inuu5vCLkDmLJHQWDLEBexob04l+8ElqN2K2R+ATE9QiPGXygUxNv1WV1pYy
gWG+17pkINPoU+fkOLeDZa6salUm4qZahh8ZkcwHgEf88QIhp+M+Oc7IUqK3QO1q
z0FcI37TstcpXn0AHumIlfy9cXLmlaKITHDr8aj6V5n9761ppMZH83aC/igKW7xm
frt+8MyQhQKXPv8r3sC+sVUbJvMyRstxhIMz0+R1vk4Dz4Ypr2itq7ccKnaQtm4j
qqqUmfgJ1iWW9oKXH3rz3lxqDvFKfUHnSJRZfEqsI0QBQSdHZyMLJno2WYeStyh+
sU4WwkOyFbZDUQs82h4LwREbhQL4zlmnm1zTHn4/uPV1AlT1TS932TX/WG4ZVt0z
XSvMTzvqq3p+HKEb/K3naL8BxTZ/qyTar21supz/LbBj2ODRRAcgBaHzlZJPBmEz
K4uzlc1ee93KmQ5HAHLrLa2QXGmcLnFX8sOaizwPucl5ivzHufesk1iWJo4RB9If
072OLPmlIqUQu+zt4dyD38rX2ZxL2vXihS8m2NuenWIbuHV5c3eOBT4zkMv8ngAg
38v4+ISjWAs91PQalTJpAQEQhJL1+Xs1todTmQu5O2DLMa2wQ0ekLuj7rVZ3Aapb
uSkTLglUo5c+4rg8psSJKWrFBxZNU7Yaenc0F2r7UWMoxqVKcMLwtuYm+bqBNCwH
n9/Br+BqiAWKC1dHyhZ84BnhGAYCk587XmJMLvMkgwAef4/OaZ+jj75Je6eX2GLD
DhUZccx6xNzTYwpdEJrD/Tivnr+D9Xo47ilfYNMwFqLkgySoNmFLhO4zjM3/dzUJ
YoAB/YjGlyOsyr/gF3oBsyUfPu04MOlichRQImnG2eWZkgR9KHpQ2tMHg/hcv0K2
/NdFbQtYWJ4kmF9hYBrIZVMcmB2ucka5VH5UmMElrS8pMj63Il+ojP/G+JNYQEJM
xVZ6446xLupfaW937y7JAmAfemfY10lzF/DShBhpnUho1po1YhmmSuF63/i8JGvH
ZW1JiFIuEThsWlQTjGJ/D09PybEXh8xk5lID9xD/rpuncZzOmUx+ONR/GSSuXQi2
HaThr67QMPEfs9oy3+rKW9P++v9zwkeHSzUKADFx2Im2X/ZzhReJ6ovqRfs0h9Gt
Hy2/gp83ljE6dffryxOgxBiaJ/QKdnbwq57o5FcUPRxp7GKcunqw6VfT9heny1mT
wKyY5fKvsZjFEF6Zxuzyzbe2tenK/R2dzCrapeL5bwj7gM5f2UTwAeW9+/jdgCjY
JByrERUkfKnhroWM3svZXL56UZX6vlMsx8aYVxvtkUCxmnCuf1IH8KgT+dJujEWe
HcvD4g7lz+K0dwH81XcW/jFLC68X8tj/pWeC+kSeCLuNaQwo2041dt+zltF3XkiA
2miT4mDAbacw/qIXgtPkPQpJJEiUz6boUir2pPUQppstQ/xWzkzqAmtaLXtFzvws
NOwpHed0j3eYRhcRvyWbNmgHDTNimzf2glvFb3Cz/a7wZxUdYadAoO8qbmzq594h
LXEZrbtdLQVdOBY2wZOHTwNkuNwobKjajiKb0sry8sAhAUjEhQ6H0HsT6guVkvIG
X0mhNlfE0VCw6z6tRIelO1nlNOy3Hz2BukvGvnFd2fOrTMnHFZJAMyg015+kixib
tYdsQhcCrNxddEcJl+ubgnSxeHhMwh7kaR8E378oKp4c1PFLabMAZ3VlIOFPlMfi
4JyhcFY2ZzOWf0zdqa2Ej1WebbO5312WOSgtPWQLuqv0/lmEHZ5H9tNsiZf0IILj
VA5FA05OH5fAgBgEHegP9EVeSGR48Z7fU7UUZ7DaJ6roj3XZ8m9qYUpEbX1L+r9e
Jgjwz/XcAkX79Uwk4dI/Fxj+FNRJ0zKgQgug7VUAoC08vpRgbEqhrWATW166ouuS
v8vXVL6F4uXkbrbRGO9LeYcVWOriEwpRIZ9rjYdtS7KHojDKO+Api3h1WM6NDTxX
O6FvymrD4UX0gF9eoxxsevp3cZwyyHRxQxWowQSm7f2UEUCjnueJnJ7N9k5i2P0N
J0adMYBe0CbsXv+JLIW+nrASVfA0XG02nXtPbKT7VqqHDJR4T4Ee1wc0N4E7hc8U
F5YUARZ46RHDy5bwXevlPivM+gIUNRYrwCzrFnkHoCzcrJ8w0sal3oo5LPrkilMB
x2o8gKr7z4+TWYMBiOmvT49F0K5tzEPUQp2xkQOdgSPESV7TIm64RSgIpCbQbgDt
EAaadQPSAMwFgF0exKaPJriT41Su/a9h+YN6Y74CiSzmNnqkNGLLu/6Ko13Mc8bC
ziDfGlXaVXwA2s7SqHPSzRxfsi8XuVXpnYRcLBjgqOJNGOf/rL1evGELZr8AU/56
hjcq1bhZ2EUIWoe9SWE7l3W7y/K3tbTGe8fb6m49XTNUno8BpP2bif/PA479fTNN
yhD+RqDCtGFcqX0pd1J0CjvhFK6vMS19s5BQrum+Oa8gxb7rWqzraOhLQKIcIwlm
BICGWNTPz/Ct6mUZodfWXQlW9H4ytTKcW4VfmS5fAdp2rpBVdX3NPejCEVlMkGKH
Ec3XlglI+/L3xA7tvxAms1kBnGShWN8QgN044pufzKWxd0ZpvgFGZwSqbHSAtCh4
dITEDzN3EQ6PkY8qQtlfQC6u4Db/6QhXlU075ciASY3k/h9B3hzUO3mubHB56Yyw
B3kd0hUeqCklFo5sR76pP7sq5aXntoy4yJFQ3jkerz+LB7QpGqh3G8XVHWBVOr0g
BTeFnNm2LrHJYF9EixeQ2+BzVj9IoZpBrka5Y8z9UPUnRUdDHD0qRwWEegtaD0bi
c1Sk4oS0mqj55c3U10Oj64iduxRp44JJPY3cSaJTlrCPZKfEBhtPActE1uV/+wKM
UWqpTe573u9XxNsGf1t+tI3//7ZTEu5yPEOJi1byjmQ+ZmWOy5KVi5qB8lLNauEB
dClTbZkSztvgoD3+IhVYX0CiCjja+kXhCvBimNYO1SH/zlDppMsBEcY3+3nyeZ+8
LOSEpzuRy+9rgdocY4ynrFPTPgtetS0jiFeA0Y2HUA/sZTPnkPZRk74sRSSIRKzC
ZDRf3yGTC379/0WO7DOmio40MAe4xVixnweuE1qsekqOZhfQy/jNlHcmveSoe4EG
LtTtZaGF4/bfjfjXvw3OJXzKUNP+pEakwqvLfW4p1NkovSFTda/Sgur81Ezby6S0
WQYjVddHhi2x0saw9Qw6BB5T/cxh7iLcFdOuBE22UAOQptmXV19NSduzr3ZGHegV
GXwgbMgJakmZRN9yk65XQRylwe3nYfrqefT6j4bJfpy4rmKMvEO0YXgEVwYX5/QQ
zSPwe0TOg41Wgor/1YCFC4ZHlZWRyU5ibq0HMS3dy5Kgst2mr6nYdAF620zxg25z
5vRiVwrCPXCHtYr4wPdXnTQxeVhLWl5Y9zzcH4TADp66XQWLtaRirLK/bQoSkqIk
D5JsX+RLZxgkwEz1m1ycBr/pekoi6NKaxY3U00JbjARqn8aeUwV9lj7vMkUhB4LZ
PWwzyztdeyQ70Cbl/YTtY2/ZY72QIQMO0DAR4Khr+b3/Ix2ViCVSj7uW3jJnG657
XXtuKSoeCWn8XsdmK167lcZBUDECfTlwFABILvRp7U+3bs8z4JfbvyDqMv3c4B++
oxiJ8VdcESz42GO6ozuKidA87Vrpq1HKJlxkCnpV9AH4p4M6d0oW6xT3jqzPK/wC
j4zte83VeUbajssLSX3sjny4QPbu4L9JFqo6g961wRnt6RCOkXPnnfQE1GNhWUGt
iglV+M5/Oqgjewy4KqZqgTOfGo3hOYpvkDMtk47i3pqy5oVSr1i5ZML1FBfIMwQi
q7+yw0r9rvpSPF/nyPsvEDoIgwEWuJt+GQep63tvmAh2xavjEqdMBhaG7Po7R2bg
s/Hzsm8IwM0QmYG11r8L4ZUZmyUEwpDQ8usujPNehK+6VzAdQfCXexJigphF7AEH
p7Q1qCrvhQBQaOncWYUAjxGBKeRL9AKWJkC249kkunh150jSckoSIxGxYwB6pWSR
CUaXSzgp+GowpeyQEyKzRzKOn4dbI/5vYlCbvgjO9RigbKM0v/uzJ5cC8DaeNI0D
Dj15cIFeHfZ7Ka0U8KFoQYA0/q9ltnxJMRfPUyIXfgeF/X4et3wKdBr4fljFCh1f
N8HSGSoU2khCTXQ+ofS6MCZCOENxIpwsPpFIIYDmcxk4JLp3L4gh47zcqo2J5qJx
k3DWRBnkGhzXHy7pssxQSHdDWw7l8SAO2sbc6ZVFjorKEmCmTX74fWVuJ7V5UeLh
L9vCPiS43Gz72Jf7ZcKaSDejxcN2LPGu6KTZ+A911qbDuXEwMDoW382Xkn2Wy2EG
xb9/zMoI03cwbOyzZ0ltOejJ5WbMzKh8GSwGAcm3S3M4h/9T8iET+ikBDtXU3osb
MdRkKybg2lZGpJ14VW4NPU/NjcP96f6ubo5xYkvC85S0/IpvwcCZEOFGA8WBsFNM
W1glxApSnKzD08TMxqweWQHw+315VrHjceNA0UhP5D92CD6tGxbla77Zz7gQnbzU
qQasWEoGi+W+g0BxSnF5wvG0FJLUPtqzSGRJkFBF/T3rf05HLwthNPxNy/fAuLG6
u0vIXL/Xzh9UMDpB7S7TNLvijm9rVxkfPc9TOF/OSqRsjVogWCiNin/IiAPaHO04
qXa/Q4le1Zq1C9AT20exm/JJ6SfEn2NcAYUnIby0UsKzNZ+0BA5GFzD2IFQ6QYkE
YUPxpocbWEzOiDQ7QQDwDj447ymjNDg7jXwdk692ZbrYcIgs8F04qpNq98mOhCM+
gRSuOTv2kd/aSUudC6d/tKnZVz5TURFIyqIzdF5aQ/RODyR+nhVmZ/5AmK/9uitD
jfGEPTHKMMphB4gbpTmneBAIUdFy1YVLa2e5yTga1k96wZIVY2CGeogJfMMI++01
VUaX5ImARByTCT8qdSEpQERUKr8aNpahZ5Y6KhhxWK5lx/YihEX5bVnzcgfmnnT2
qQOyWKzjZxlKgzAi0FBVJq0aaA0aXnniC68WlV2b3XGon+Fh+Xj3rN0uObEdSjVM
0wRLV23/pq/oo/nyAp87mHjfcji47dOmF2dj5KI3ZCwJuft0DO+wR2TZ25oPLKD8
159ls/eZ4lYo9yah8sKsMIyssXvNytxb2P3Xs/skqEqLgFUnpzgpv/wq/WGmGLXH
MGypYUKTYm4T1pqfspmDgeBKijQcxdhel9s6YR2Jgydg8YAbDkgj8IrRCXnUPGxt
qwO6OjJy8L3dYQckAZc0r8csj66DK2pV/+fdlxODD8nlRnmRe5nKcI1kEDAyf8th
XW4A6CkQbozxD7Q9Z3bKM6i50vXgbNzIfBp6yAXj9Vn4XHuPtXGt5xP0dp5Wm3zi
VYigLUMiFnaeMj1qJhbh8UXMxerLFRE1YU/0CF7MYjZbEirJnxxt79T5/mv4st54
l4Vcw7NEfPR/3pUQzuDQxpvm2Veq0LR1PD3so6j5WMVMAxKNW5z8ogbNhEmQx6Cc
wlluVAMc4P0eILn2MKzvuu2Y0NQgbU14E38rvY4YQURrU1RiVXpbhJ14zdg0ONrC
oH+qem7QXl+3dqXbw78fRoZ+9Nv0gqfs3zWB8ce9IQPIaQ2aC5LShsDL33cJ4hnU
fkdIXvnMB7a4gcsnh2sab04fCrCFMoJk6I+KzOlOs+WwIozihjWaERwBs2KpDave
HML3U8iWob/PHRQ+gXtpY4XemazJPbFSF/eyOqNjDjPsbU5jbjkBtO1/6w6nqh29
bQ2i0Gbi8qKPiG6fYZF0ZIF9qLRMp1SJTgi+41f2e6Er2P1Z0s60kQUhsat7JB8k
tN7z+9Cn40GWxUm7sjcBHKeJehBhvnhMpNWIQwC7NuBsS5FELW/BFP2t+AgC5or7
sL1fgmrN0Z+wa+9RbRl9ezip59djSAO8YHoYPOOepwNpk5J9a559FKvw0OqXUTLw
5zv0XstziVgznQVzmlqCwMi2HOS1DgiMdJHMDZYn8TpdP+/gP8+8oYe1ba21fZ6f
m/9WKuwrL5n9NQ8winWkEEk/E74E2heuGUrOpF8YdJt5ofRhvRJvFK+onsD7DvJW
jLN6eBhgkOus2plc/ouG7/wgg0AgcnmdvauBheIwTSo4gr0V7UWoNBOM2raGO5Dp
HvQ27IKn29eMiIcwk7bPYDBKLBLTMdKb8EL0DVhGB4klTKjVKVVuQnj3U8Y1eIUd
FMvnu+opqdwOUOgPF9qoHA0TP3s49JfCGSFOjvUS2kedmklzqHs8c8yg10mwxNSM
e9ZDSrpBHsXFNfSYYiz/EcI5wn8It9sGCPIj1zrj8+LANM0Y4UD6MBFikhnxCDES
pgfCDHgLXlsW08IyV+B/jqLNbvIaplQ2bNPGuQKa0UwrU30ZMxTDzjREoxrUwZ8a
h2HAxNc9x6OgIBeoG3ewME+hC3fQC9fbe5ZiPP1r3057oKT1y7eP9fKDi+IeXzpF
FOCdnf0qW1ava35o24st5WPoRL7fV4Tv7FkPIZiNDh9z3doi7KsbR1+fqYbKeDlv
nStnfRCzzVfCW+Ia+YoFIM7W6WFGHH0N1NAvMZ0NZg7neQ2mCSVHe1UIwWrerJxK
41wG4u8+yJ0dfbpuQSkqnho0FAkkaNw2HHKB+FCDwCKiFvBSfkSEc5wGP0+RNF4l
lgFW5fEP8XEZyRTQ4INUWU9x9HwgBCfcvhnDPTpCbvD1S7G5zaTCRK9BdMac/2fs
5RT3kjTNHFmhh+EM42F+4eof19x88kseWzngMR+xVsU0CAv7q0352gQm1s3Y+NP2
iHasYXc9/1uKfK28owTHZO1FfuZLsrB4LYSM6CK2Dtb3RfQzT121weRMEkOgre6X
V7dpp+GaWkHmPdKNBrS6beXS9Co8qhKS8QiBO643UXR17LIcyJvrO7mgAkvcdNgA
FbPJkWArZZrzaavlPIgT5RntP9zLeWTjat+JgodxomSIHWIv9AuyLe2NLiLUQFNA
nhR0sWsOEA3UVcxww9Y2FJvTZJ3LUTu3M8gT7uC15QRLrAAuf5d3VJg5DuvVamaO
xs0CxLe1oEVnyj6HQCNvpxMrJt5QxznohgLI4iyJXgEWMliG9ft253zkTAzv/p4I
Xiwz439CZvEeZizbRlmMES2dFoB3YNnjWwguLjUaWWCWivotP23J5vfpJkKYPePY
cmQDM6CwzOV+yCYd9BiS0CU+aNObEQfx/egvBDsv9Fek4OhlU3N8SHW571oUE4Lp
MCOpjs27qdzQEMUYnYfK18e09et6G5pV/VCIDrBN/XBXDuXcFpeTFYBeCviUztWh
AR5uB9uwGi28EzNjvDf76vkNhJjE3LdZrdqUx1Bi7fbXd1n5lg3Oc+pTQkFC/1x0
iW9I+mV7gWmYshee+BhFgHoTj/3A/9npStT+lkdi8gNtigc8WraMicLCQcLhvqAz
kPOICsncjbS6zCZZmzH8IkI7eVHPSUbyYIWKcEf0T4B00I4fBwhc8W7aw2z2YfLH
zBhkMHPOYN4lsyM9Z3BRqigZKakoxNbMVDtk0B0tgKPQZ1K4mKCEuvxdcMAq9lqt
5m8x9lH+8TiNXGLvBW/IP86rL5WM5kEgDKhHllOoBZbe2oXEbOu8YyklaR3HSOHn
cV06sjcNFGLpXW/Eg2/Lt3ZE3jbchO75ZGsMGIosopMMCfg2OCGNQFSjXeuarqtR
5cxtwJTBw3w0pfWk1+9VzJcAawnUtXYFZWjJmNQTSNbAob4la+kEF8iq3mTkDgoN
Ym6by9yvnhLQWnH7DBF/yu9mxpzbM1+oiix/AcQE0Qo/59xqeDVheAswtrrpCymn
D6QTv05drXWtWvTbdQetkRfY/KZIkNfY2xik4py7caa3OacJw4+TWx3QTlRVaYul
kP4FPkvKSCYm5ucoEvyb9VRS5YMZSNijKeYlZCoPwi9B+ZSC9KBlLCzz7ZJ+JYfB
MjKf8kdMFhLyYQtpMOVdGhToX71puw+Czxns4zR1heDOO7wWAWBghtPiA6EA+XdA
DZ87o9qp/r6tn6kj/dQ7vzMj7kBf3UnNedN/Rl53OESirxnj+xhsY+W79JVHx9Rk
Ebhvx06MylcPhhuBTh16kskv5yKVaWhXO99vRgJ8avvk0kGClgqpWPaUmlWzH03y
c2dyxEXpjLn86/86wTHa32TH+0gkap5H+ptkEsWvgY+zd+brsFMDqARaLQYiLVir
+05ALMu44KbgbGDo2L0hxcY88lK+BxKkIg/g2Oi67LjWbfkUwk2N+Z4OV/alVgM5
hy2/NENpmKyXg8sfryhkHuDRRplJS2sDoZqUqkNFSbL7Iaz6O/A+VtLMwcm2kjYq
cdv+gN1vJaWpwNrb8InsHPidcG+Do8Dvbuw3XC/iGoxobZ7AhABiJg/GDYoxq5uF
dHUWHZC2H7s8GncItHGRFKT4ZLqnj43SCjRe7wYbchvQECLdF1ZXgdv0/+T49WBL
Cg8K8yjy7kdCmI3Y2xuuCKjH5su1bqTzDT9nnfHD2Va9ffiyhc2vbED5SW/SBZZH
riLzFNkBZ65sHJwovAIHQjis+Bg0iPZp30MhIQdzOsZHPGUIk2bbpU+CLndTrf3x
oEg2lFDVKWzsBU8By7xsec8J+Ohu4oaE6PnWwu2AdMwLc5Axf6VKFSQ4cdvlqnhC
nIBIygKRBZAAxWgGxaNM+mjB48nVW1au5UavcVu7IitqI/iJkbW3RP3bOBb788B8
fRwZ/rLN7bBP79HGUj9I1BJRqjj2nvNWgVbVsW4cVYGBN8zNrzZZ4MS+218v0ERQ
j80dl8S/ajtC/2esfli5MTOT/dVjxVxXPo9mU0jrTj9MN1HLyAVYPmc9iZuEn7pc
mmtmWjrOrsEWfsJ+Z+k8pz4iNRuVrbH25QTpvsvpwNlMacW3x5mYkDBJpFNXagOY
VdbsFDuMombarny72B4tZKhR0Y6JQfWyv2ddZGatJ1vbM1I0CF0XDMW/u2lPq6IX
91hTWP+TGQori5iYdOFriKq6YrKFW+zX6jzQA2c5P1fBUm00vL9at6FYPqumzVMy
ogS/4v8o5ckSzcQ7W120/ygIR+wwSqmbcgk1PtI/6uxkRc8s97gXsyTEIr2Kocuf
OqiYIem755FJOxBFQB4VhL1mupjzZWLmV7QPW+Qi6jx1huB9WVah4eP4GazeZ56G
YfadSjqJHJc2pvYSNyKnfdU1+jIpsahOCaZajFFvTfUyzHFvQhJbXV1XWaiNH6ck
avBgTORcwvxrY2pPFLQQZvYam3+VonqTAsXUHXe/S6lRQYmIkv34wEo96sSM8KBe
oU7hA5PDQyXpOgfDZ9qf1vpy9XpG+4MOjpy9O8Dk8ftxchkVwn8QIPZlBz1M12oU
RUAdzv7crvp0E/oiYgax3xsQu8zyTYd8doP9//4w/jVRmEdqo7IrBJtutwURtvat
G1DyFO2Usq3yivYduH3EL8VqwzUFcCogs6qGvBezUWL+aKHs2w0iceTObe5BIl4F
rPwCold/ylfteJww/Rwq9jrlLxcPlTiWBJm2ABHvQMv5R3hitSt87bM53msG+rWF
f7lnRgjTT0j2/8uTPl/fGxhPRb7fzoWj2I0X8v+v4S2Ijne67tmWx877RmbIYVCF
6yS4FFuFhtmVYK/kdbTZE+iLsICIKZFMZGsfdnP9GV0rtY/THFMj2dFsZNxzBDlt
I0Ars2D5e6DxjtZAjnU39p8g0Q6IOMALUuD+72M/Aug9Bi5wCMv3HmYbEmfa0uJ+
4Z6v9SGhZFrMLzePHT9R3cD85wLKirME/rRD9jhmC3KvVVKMI0jYrDx0JO3TnCcy
dtu2nW884cYLmastPX7xFTaFKl+OYnVHRo1Lowa2Hp/rOMzAMQajDe1lClRvDRz6
/SnVIhpVqmg+XKkH7F+m/PUoj4L210abFNjX0HewcZZSDK4poMCxw8OcpKGZaMyy
0zyQYA51MPS2TugMoJFfInTB9Fpt2AXFmQYnDSWCVzfw0U1hovLjTosh7Knl3L0B
OXPPgK5cXCExvg9lJOTKAa8nbOqZStya/BsO8CtGGcYlnKIudBEWDqvFyKQl3MlC
rSSbj/LXLPxclqR/3aAoqF9tFJ9uifC9bWk0F92Gfqb4lwAbdztke55WQ4Ussc0I
OP31rS72ZOkOMXsfx/0BxUMyPeZdfGkxJ2QurrjevsBAVKLDLTT5pA8Wo5yUmtTi
qyje/jEkS02V0A+lGadug5KfD+QIuncnSCjLZE1b/8bYavYP/kjQrke2qqKfJSQK
9koX4MXurylHHwz85nQuUrw3IKxS8xiROzPk7LtjxSzvu6ZDKrzVo5gyrGteLRCS
CbVPVu2rtPxkUy1W8OGM2Efqq62PSEqoO1pzgSL5OpuJ+6o+Pm35+BodfOKkfrNi
kClTtJGqKigyahqgBAMbeHssVkaGspgwsWe4OvzUZJCoVPUJT+FNouRcvyoZBcfS
ix3vsj3KRw0wSm0yACrzlD2eqYEgQQz5+nZshNYUv+Ubjp3KDM+hEehK6CSKYUJj
dUIW5TPwkFTJRumXELon0RhLyG6sD+64k7rkTSUskURYtgRpBPYq98tlV1lUp79l
/R4hapKbOGfIu7FxvGYoCdELTuwvMjeLqM0owyzwqT44JC0pauGbJ/LgDikIWBEF
UMXwLkqS/9zCWHTJsbTZmA5GqeDeI26aVuOafxCl4eaFisBrzWY+x3p+gW2+LwXN
pAwpQ+StxpYnnKhZX6qAgfavWEq2rPEcEhGJc8d7vGYCV+hkrDa7CwYaJOIrOuh/
q7r4YY0CqRFhDplO8aPrLlBhgOm9tJ4TMmYu5TTJV3t3ic1pkDvZV3Gyj7zZ163t
XJFHx0S5K+BvtD/ENz1NrpIj5Mfg6Q14oSpT55MHvusp3nb6oCRdAgwj2JCcZdpY
I5zLFP9e22jvjql46D/I+CH3nB9GwaNmC0OpFxSDkY8xvMOi2wzQ4pRQyf485DqN
a8zuRvFV0teu5ZOBZiQR7xJCvr/zwU8BxZpxO73nwdQbSxIf7N4ES5Tahfvb9Mt0
Gw/d72Oup+0f+8ujiFKV/dt53T96tw2k/e3yZ8Fo8cgGalhYm1BWtkTftpkvbczO
aSDYNyVtJth4nwIXZRP4Rrxw8mRAbi+LIHn4Hf3Aqi/xOYZgxSIrSHpB/38dHCUq
KLL/ZaHDRZH2OmOjbanzKQoJCbJJ2dGIs4R6MjWcJTANOOUk6vT0x6vbcv/eolnW
L16iBDUCQ1o93KTza5JODUNsgx2N503FYTK7TEtp8wanK3SPiSp/1aQM3/kylX0v
N+X3/fKsUCsnZyYmoRjVvFR9+1bFaE3ixeCr0tNB87wEO7FQDgUH9qyus+sql6pI
4JuS2fYcLHEKgeJqllyaS+pz1+zSPQ05CLeH7dIkQlCdSeKB+2q+BTLgCP1Jc79r
DvhbopIbRI1aipseVaAVbPwa3NqUiPhSZdCP2EvKZmcu4FERoa7n34aqPsFrq0j+
nJpW8DItWGgl3Gza4Lf1K7VPODEYDo5okzZHlXhucp659N96h72JfhANyfvFHCqU
glIbeCpKSJ5yRr5V95ncHd8mWK/ZefVQ6hYO5CLY/oMXCBrOLrK5E0NzTMEdgtIS
cYL2HUgResnG5Ul7f0qlYDQoKMAnwNeUihz6j1BF67kSc7XG1KU45+yY8MR+Mgkp
GwmAWl5LGVwsT/emu2yecaUoB1gIByROMwDjrbhMjYl5jQJ4O9uv7GqAa7u3w80k
4SbnWuov3XKoNnUixrUwH/QxiE3YOarRxw63HjaD7BkhvvPNKBK9p+sv4CkIkbVx
wY4byXf7LM/aTkLwxQocFfpfxVJFSLcUVIVAXmbxrd7wZZjG9KoTezJgdX18p9IV
a3jUNyHsaIHHNkTa+NNRgWhYm+qsZz9c397Arec1+LOhtJ9hflrlnT55ilAgYJTx
ubB9n6x+n8HPKhVCnYtudZkyJCgWBTuV240IWQwYWBFFtg2F4KNHir8zWMD2xhy2
jnK0XjKkj5zD17MeZa0jBDk3jOYtSohUBjlnpwW1oYUt8gd7XyP0kImiT/RtjoS/
yMjhmd9HvcC6Qh0DySq+BLXtzo1wShM5hVYhwUKYCBLmhgmqE31bcx4pfa+VwyRf
pF0lCb0MMgwJlrhKi82SwHf/QCXpc6Za7WBLeGk2w8NEYQzsyLP1LvMt0M34dY0X
Q/WhwSpb8JNXMM8Pzp9MQIYStomhlMhFeMca0gsgfjNFH2iIej+73zqbPrSaJUqh
QgqHu5iJENrJqIjoAgyoVmUpLeZhCjeFoLBd0d+jVJG4k26eMwbxWDSDckgxQVqR
4zb7AAmVefhu5HaSqfJDY9xXg4DdYIhZEoAJBFOrqZjP5nYhVcfZmss00AzuO5CU
jFe/xPSOcrngerYnATQ6wsMJ2bl/EbGEINx5ubfvddXpATickHg9SDsfyNoZP3HN
EC8iL9WTOc8xW/BuyjB3J6oamk2ok4Ac2pfsqrfSv9hCGgad4r26UaPTRZ/j1C89
9kyvmoz4PFK2J+2UY+gHjdJ4+tQa4tiih3WL/8/UDjSY2EgWT3vhE+GR6nxCWKuE
eatmmF+cwFjg+i+6ULGQgGbijWzQOuCequVYsXfB6Ol0enVHvsCwczBchRemNIzg
XJPRYPngal7+hvoKW+TUsC6ygOzBjCKBVIH7RfjTZcnvwf/UW6Sb+62JfPwLwGL3
EranMzAwFtOJO4gisACKjmvk22FuiRysCmsx/+61MEhcSiXzJKTRCBaFYezwuTXD
y88bpee1ejNuHyFPpt1VXRnfh5/zyZw0I6Iw7K9i1luHWcZNvVIUcDYwQbnqjz+2
AhKHm8HHP9B1Hk1GQrAbq1nKAKMnl+MEQ4K7MLKZv912Sk5liiARgpp9G6L7khOp
I5Xv+efsBHjEEEQox1I49p+v2sxWI4125O2GN9xkCoFLDsWl/NcJWYvYjhC2j00c
7t3wBesmiZ4SR3jzJGqbTx20PCRAFOJg9XRKMIrrKadAV6lMqnRayQVuDB9yTrTN
PyFgkIVjPM9zad3cPQPKAhuftlJWLwjOCDBNs4XRwF6THOFj62KnwKiNbOY6asla
O5l7s6k6UsbTQpnJzLn+galKTGYVW83J+Ib4BDgxzQDRnXaCjEvUElQP93j1cyVR
xYyKZlq85VSuvzqXJJxvoK/eSmTmknhH9EgVuYvzVWWjMwviptyo8LE5crgtwFCG
jdcfX4keDCkqwPFifV8qCPLOBL8IINSXOf9vIChsIXBSeUWGqvJ+C4Ocb3H+FFxN
9Fj9d/kJVl2JMlFM6BNDczne1H62BSVUgB59AVKaNba9aQcLS/d/gpNGYUJaEx8t
6WAMov5CLQrcoh94YEDkZc2Mx8LEXoS7JRy7SQnWdihJ7F908bmWoZM8Ou3By127
AsicqcOM9hgL7rMSMAvyGcyBEdFUHqpfIxRhiNxWYX4Uda+d7W7JWgHkHgivkGEv
kK8PeDorkzyt2NVanGzzYRZ/Lj8/rRx/Rv/CwL6WQBnB7B9xs/VmH9h9t5Wd6SE3
YQoCvDELBcCYFNLmRZqZK0Zb9sbg5tk4oVQ/p1b25IUi6jcMrzN9CjT71hdPni/V
C9BdaV25QX0J1HgE9diLanqPtPZ3BIgsoMcC5L93S/VEX4xMea4LRe48APLkMEbx
KFpgqs7m6q/zV4m8YasBMKuhl5lcOsUOEfEJYDwB4PAJZM1yc4xHimw2G5knRVmh
fLJA5AXA/7bUymgNNYRkk4/KiCFX2WyKnHulBBZsj76ExE0OjxYeL9BuTJA+xFZg
XeWv4XG2p7uPSujqb0EUuIhQ7KwZDCkaNtlX9bJuvi2N/OJvmLRFMc53MRz2nLla
yglKcpENVCHf3XkcYuKEZTRFdxV0fp5W3R4XR5ChnaXzdcHR2ADeCVkF5BHruMVJ
nEpLWuIGN2rFGx1FZ065yKiVQvH3SimfwbqMcYgHSJM19xVLfai9zTLN8mGIP8ML
K0VJdeHDiemvb70kiYZ8jBrXxqgC3+ZkkxoBYxUQFxKSKiZlh8qiAqVUWOQIDkeT
bMOl8nLKm6PDnm1VZQg+7cInlRuUAWkO79VBsclenRyU+0D9ci27IJgzwfBqyrM8
hEk8It9DSbu/ZqiDtJ49jUvziV8ePppad8r6X356O3FygZWOkQkAxS3jItNTBhDu
FVAstNUMpAe4bu5dggC4Iv0idDGnG1Ssrnnu4EC5zvo02gaLSy6dH1DXD3CGn0eu
14wLXBGY0MUJ2jH+qStFk3u8NxxjZa1t4GZlxuUQ2xA8Bu21jHQ9wD7sDtd3LHit
OM89UtN/UvI5iM5O1zqnxW+OPh5pkW+iLks6/onzVhK5Hf5PwVW20da/4V8cP3Ge
LKFcbm1cI35wIzC7lxMTnrUICuL7Veo9CdziQti6Tpla/b3BQCZbJf5q8HDRshgJ
g2nRHXV5oqwjxDYrQv9Q3wKgoOdH/44NeQy4m/SRyRZ0O6WRkqyaf1J3xA/5W5f9
GGLozfywVKDicWdIfxGujhBUbnGyDz6HNhkfYpkX7/9LhW/h6gHU1G0QefRW3Fea
Puj+oDXLfQPDjncjvkmSEz7nsodd+YHcBLBRlftJrz5I9/PsvPTgQZa/rVJvX+Ry
h4yC9tsXdu/EpjYw0TReMhLz6VJ32p9XZkpqxv92d+9M6xx5cFNkGCdg8BONUhiD
jLadXRn4Ypef86iGuBWK95gJa8Kw4tbbDI2nJ2JnrgwRwr6E4TniwSRv/FLuLIcA
7lJcZ10kBaCsjIL/HTUDgQQcoG/8GY03F7FMW/i+nO5HSCczSOpsN4mGUqTrtrmp
OV278mOFyz6YAdG/iBg53CReqtLpeW4ivWBOYfVFI64Or2LhCw1yI5nHCbajpNov
0ViJqLfpILHi7tZdRmIJ8VfMU+N+347Zs5KxIONzZHMhK0xc2ZSUXnfXw5R7wyM5
eiVoPfKDe/Ie16HWnPcoeQBw0Aw9x1h62zmzx8xzYZNMnD0EBnsSu6wGUpqgPLcv
I3F+x12xgM/LDVkk2o02NJEzByHvoNzo1pxWsztz0TpDeLxpNcdKS9n0gHkv06h+
`pragma protect end_protected
