// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:01 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hkL7h82TiSp8ceMPZoR8Q1Z84CGVhHaiM9PDlJxXEYJIO6SLH6SyPPAHMFvvn55F
9A8JvvWMnr4/4Vrp3/g2r409VAimTrjvqSG1L+aYSgRpKozpex8B/s2m0oN2d5cx
MO/0wuOphKjAKohkeLum3LCcAkBkxeUaJCpcE0MnV7I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30128)
1g8RwRkVjgk0ykK3Ktq6bq+ZTvC0P9OzNJwgCp6Ijueb/BxjvR/ZF+3Z8rjUN/KO
vfOWpvn6i41PU5fW+1RWYt3CX/6mttc6nnZ2t8yVg/PyyWKf0V9HYHw+BGWtgUE1
sOHASIaOqOWBynLXwYyAcnXPKvlV0yOrzccmqFyTSZW4eyOfrFgkIAXB+w62Ocxt
VbvxJ5HVx0hFZ1DReaioqHYT6xbYqksejfEP3vZiiNkI6fTg60SoNmS32CGdvN+H
KS/g3/nv5z7LF4qcMnzrlo3bLBOHQzsKcrOctngjq01hA6nghgtBA+kugQmIivyq
5KeFODO4d0fapq5wR6RRyqOfPc0uF8BazEpor0gDek3rWBGKlj6Mx3nFYLinXWGk
ViB5Zoij0nJIGZRVVhE1DrEdM/iQ0LPFfbYZJEmWbme8/t3yx+orOhquOdzZBS0Q
kUX48pb8B02nYuACRIWofQCzrA9h3wGpZDu6J9S2TkxDA/B0ZNoj22pBhHAIxFnt
E1VmykigUeMvQCz1XHvcvDeM9cFkj9mRjXA/Bk6TEWePrVRLh9VoTXkNxzmDX9g0
vq9173+OAw87RUDUanhYONpXq+m/qGC7sNhN7uKiDw88dSK+qCmFPxY6s3cHbYur
xlRmbPRpApWllLYM05+U9uc61qRlnP6IUYku8mgzwryOFTEacjgIDGFtkrBHLkXP
Ppr0e0CZwdDJomoN/JvDpIyBPxxDWxC+FE0wdSkNweZ/YwseGS0FeVEa1PcVjDGk
xPHYeZ89Gi9/zKilvGTA47t68jyWeW5/r/ABRdf2wMrqeBja7zHMAOZeFzFbyT3A
mIEMNFWk1XyiAxyieXifGmtUQ+fNdK62dQfbzJAFrw7oioG2iWQQymc1xlhFV2vP
Pm2sWBWmVrTLtAN6QzExpIMHwQkaePDK8feAS7aVdL6TaccaTb/jO9Q7UTJLv0Rg
3/aF67R3X5kM2l1yCrRK/Rp3SsHiVZBWUJlT7MPs1i5b+ghqBFUdyKGGXD5D78f/
r57EHLPlBnDKMRteUOaA7bKNqX599I2UJGkQ8xyzOQmuBU/O769ECVmmblcpTJ1s
OUFCQauGKOvHq3l/+xq2UNVkA84Wuh4XfqiTYNLBYzF8nhK5+jB5R6SrGTLosW1z
KBB1DL9A4W2LaooUPaDxDl/lBuB3GU1n9J7spTksRQm5tloL20ZTPhbFx1hZ5VcI
Jjc7lcBXoL+a/EMDAj/CNX3rpFX6Znhb9l4CFudS8R6lvO85y7dXPlt2cApKuMId
R7GPcVNuEaYSDAczkk5C/KuDvk1vf6SLzdlushzF+AICetQKyosnqTNLB/7TpxKU
dKJovQ4UQc6SRjiTjr24eLmg4WXt0yPMikDjIRB5Un2+WRvyOBV/igDzHCiGcl0B
mGq42XwgBSEv1zfAuGoDMymexZNvXkM86N8/qRsC6ZwniAHkLkGc96QlgIneV5NG
U6iCN3xiyY3gcqEOI97UOc29jb+yMDezrl/T2+T99Jjd7vnNdyWMSM7bV2doqLEs
UOoD4OaYFTwwtsKb0QAbPCxoHL6xetZzxJaEroUxyvE4tt22ujfgqEZ5ECiE0rhm
CP3OLJxWs3TrILz1NLdO6/03NsEt+fzO0h/pX4Px4dtceum/tEAHQhwozreI1UVd
2EbbDZSppbP7lyWpJSPKz+s0C5K9NkWzPxWoc6Mb3M9WYGf0KKEjctYk/DrPw2er
xzFtbvSIZ0QFZ13TU/1mVfA/1DoxwwmpP2LzBRZt03rwMlqSbYD1x7iSBlKtO+q5
V2KrQ+kUx/RXvwwxrwmUADQio55QPFWFwVgy35YIjgl/LhB9Oulf8+YiNr8ls7ul
kaLMs2v9APWtf4iTo7ZpBaSWvr0tJf391DssygNhouA4fn5IqxDP4sDmOo/2YnKv
RdVRvjF2yYPynA3AIKSWXxIMDeukH3ZCFZV2cQB2DxUf6REPzXwzMIa3Lp650Nkl
9DP815ar2aBXlcPYPR7ceceU/WZ+uCPs3ZYVxhiUyO1WIBU0SDUwUICrhuMhESEa
P8nnRZxWsLWLkec+/PnwWqnuHHUHYzSKCQXHxS5t48jl3GefAo0iVy+Di2hDQ4tQ
5+OSf4qVXPf7cFfxLXSqRweqZSFj+kwtbVo3Kd+g6YDOOiIjbGQmuhsQXlxnLbu8
3HjsAsT2WvCJfFiWy0agBKycBVpyCVim7EAEqJfPhy/f0GYy5bR4sgFkIdjpZJ9c
DjT1EO8XqQCYaYsaYn9xN4HDPpXpRhhxclVhsSt6rucvZPRBOtPV+w5Bvc9gJYTT
UOLrMX1O5vm4dJEubMoOsVCTUkECLV106sKYXcumIv/nf33pqGDpSqr57p6YhU9G
nZpi5p2WeLke7L/1XaZ6aYaDaCEA9gCwo7GNxBMyax3uXkQoRogOg/E/SObLp3yn
vP6zFN3JQt/3UltUCKB6dzlIQphjACZrkNeGbR6TvtukHrtV9wwz4GmHLgPKwYBW
3ys+onvQo9GO5OUkFtLFKR4Zy1mMoGk5HdCmB2fTLMfi/26V7fq+jqV88DS8U3jR
g//32u1MpSJOn5tXcqidb5vfDqQL6LI9kJQf5Z6lJc0gDSV5ak0J5JIXe/iZ8ulo
cXLu2in1HdWyTcYsM59RFXjoS/PIQRWgJZRurN991zuB6ciHDNtSpRyxfMrzKshr
QjcFFNdF7Q4G4bbtMAGLJ1LunqBsKMCzbSXo9v6A4KpWdg5HSWTFbDZt/AA4fVxe
PPwthpR79U0QOEikYXzjY6tj7AD/FY1ZcfRIPouxCkN9eCem03YKHlQGhy+CUBTV
l3p+u2eqXZpqcdqE5dntQXwKw1HYD5kjH6XcbszkQUj9JO7Wvu1RZLS6bsarqUh8
lzqR7A1nZbhM+2OGdzu+M4EFHtOjy+vP8hmttIcHo1B3v/fcM9Dj4KzLf1thVgaU
UobRBLBFbP6lAC7SzDncUUNPv7zZ92DA2t3f8ksjPNlEWW6CloWRuTPnw8lgATa4
Z2z+jm3cvAKA52JJQ/tr7vlQR0HjVbyy3SjPLslT706u1NZu4HIfVvDKO33zwf//
zxdp6L8KQURF4Twq8fZzONNwg5Ujh/2eEEyzhvQEGLUww9x0pv5qlN9/W6JWGHdy
Ek7cvjD1rP8EPpty24FMTE6T7blra1DoZcxnUPbvpPxNDQt1FvXqV53OJxp+HIfJ
Nz3+E+SGONxb6ghY/Gf0ZgTqlTTjZSv8XZFhfBgfn7zh+R3sxp9pNiuVGaqe1qTY
wA4R3EgNmAhqQVpXXT7+vGwNUknBI0bD2yN3S1gLW0N4ATbKrU647h7A5KS0tZLm
eLb5Jbp7hqEPiF/CwHQ6Dt7bwwxqQiqrFDu5YzX6jeewPZ0rlV7h1fWFqkibTQaA
zvjlqnLz5rz/6sb+PGus1aSK/OTNAK9SQI8EONfzjvu8fE7bVnwICfLKZk01kbOu
WLUvlks48jYn67tJAx9sKq+XowXsqm9jhMpjHsfUqcgIjp5SZUS6GOArmSVLkY1A
qpa6PoBP/gJRJRt1nGGm5OG285xg6pAUO9MeknM4KGQxzojiaWEEU6NedPwCV67d
i2aVcrSoWS5SMipciLfMhJQ9zfgwHbsfxQfjbuDx0TOJ5G7m27qdBi7v/qkMGKwh
Mo9Mjr0y/F8JoyfdkDkWIygTnoVKATeGQC3rAKP1X7y8TylNMvOXuhk2ASBvU94e
3GtxsR7vJBlNQVh+6IwsOlp4QmmuxAWd/C+uB97FJK/SHRkYkjc3D4DptycIIAk4
CMD6KEyuu8x/Ri9AF9YH2l6Jk9kzO9vxCA/xjK5sZ/jRjivveJEYFYAk2f0o/oVy
adZSaQYAnLHRNk1K669XDQdNJMVO75Rr30L8/cclMMWuVM9wkzV/cArwqrg2ixAd
kBH6w9lHXwDljEY7jXCqtnQCjOc1LQpLATcRNLGQSHba4joDKpViOvf5/wbefdgS
QjuNbTkKWwTDUAtWGzdKfJ2/1I762PXIc5IHt2IdHCiD8ZNeMWxm5S81E1YH80VE
4vApL3R6GXIpSL2c42rYJfmVgYSEfklGRdXg/JZ0uXvAkCVRNK0ujJZUpInluetx
nw2v8dxxraLa+In1RBLlfocPJ14sQaAQ5l/3DAqjiF1ZV6iPTqdExxi8jRseNmbb
MtSVlSYu0e9x7w/P6UahFTl7dB4Sw19DvDg54vhhJcd8eaA7CSTnihMS3u9UMnYu
nRknXXI7bwu4lHXOiiIzVsOu8s7GH3gfZaSg4BYYYRV1QpDTeoJ1QQZdRqGdma6k
ePZ1X+r3PVeVgllBGvQ8tqWA9UB5BYyUnsrdgqHrF0iz+19ITDQtrGYZwgaUUrRM
Xz4XWNQ20AhNsMd0pbepDOlFqptOXYIBBbUHj8mg/fJRis1FKsfg24Z76BC9F5lp
sL5FcHat8DN690w5G9D95a3MeE+bZwTo35FChljbsB6MPfgYv0nvMKHK3b8/E5DA
Vniya+dMVay/Zywwvue2gOEmmqXS8/0/iBf6YAFGeiFinywTMHod89/hdzjNs2Yc
WR6zToz1ipbTNxbGKbiKzPH+5CbLqfNykFsHGeMkwiG0sbRHAwHw3/RpEVlsy9D7
AHdU448mLUdcXo2+Ytr6bf+Pw/J1B9je6rcbvODp4mWEVeRX9RL08IEeoD4VRLKP
3MkywtHfE45brDYzifHSQFt/4T24Nr2m27DZizGOjveXomgN+z1CPeQyUn6elo/+
QnJsaYM/xWUjTHR5QD24Y6RwKmhot9q1VNDrvA1LH19gkv6ePYMDl7BndH6LueBL
b46BZtQGGaaJhX7AhHztxyY0U4fy6hPbc9X6zFWLiCQ2rtmOdJn5AJvEWmh1PJGc
9dci17RqQV29Rjp/M61KqJGjMIU/XS08V4hDGrtEh5TiIwaZcQINamXsCmdm6RWb
YVt1O78W6+ICiuuBnx/jS8FvXhY7yAu8HJX/cO/oPCkGLdlWlXleuJ9oSMAbq3sM
DwORWPatQ2kzseu44cBmEJxjQ8+QXtwLqtcwTaot0gQFv6dbONEpNnh6el1k5uI5
bqOxOa3lfVajbCFotFd5NwHGoDw5tiJKVqRkL6tgyPHUGryypn0DkJa/r8wbRmTN
rJa9v3LzvrwzV6h+HFFhkYXDUqIxts8md9RKd6vP0x9bL8I1VwaSyKMg09rFO4mx
pTH7SMFoS5aOsWWKTs4/I58mxcDeYTcSYsVBplPa75s+hf/icAKl6RcsnnJb9ar4
eW9OY2VBlNvQXP2vGJ2FoDkb6Szeo/VA4GiopNyzpC/0UcZrksTX6Hx5lfe8plna
HipDSJqfu8m02li02JAbNp2KQtT/C+6aVlrVleq+oZxstPEB0buNZPuGFZ41BDkp
QvXGmjbDdLNx6R/ojgi5xcm0kLG3s0NoR88FF4eMJf5rteWrJ+rzntgSnx2MANU6
+IqFgjzK5+yXklHvbgQYGmlMvNA3KzsPkBOMV3pvCNWGps9FBy0ZXUgq8UKHKEKz
7dVV7hDOkehomdU67HDYu3w3yqQ3Wbg3oDj74+fJNl6X/VoZM28hmN21gtaGN+Sg
3ZKBl68G5jqtENC1lWPUuCM6NJn9B9879O4x23Sa6FYjW47t+tJhrdORlyAqRbTm
rsmAf9ARiqDFRW6I3S0liQ5cOkDtr4whUR7pYotlPupfcqUnMFkKDbocljzM1/e8
1l4Qc6ExzdIC/OOlZC7T/7YOnkMtM30s5oME2ts9c6HiBfUd8Ed1WAsjYGO8r3OR
eqTyB9MAjrxU2eqjQzdG+19sI+cY0NS/tthWzrTFoL9DdshTONmcz4EtZXlYjuXj
Ibe7nvUbr0VgLYYCjpC7L9Lv5CdNfp6BsmLSRy0w9Iq8/6hYmfy5v2g3wOWXSuPK
6+f0T1Gkf5UlDQdvPygRp46bQNp+y3Iut9K7FBhilgj/OjzMG9fna3iDL174GeZF
J1sEA5S0tB8IZFG0eiA6DIUnuT2i0VNUHR5SDY8ONKBLjygTylzHlT9ev89A8hVo
kOkpCfaIxrrx531p/blsQD4iS6CVGhLdXoViQI23WtIiLX66twJeavvWGNvTNuCu
4CCKMdjv1JUZ838+gxVSNaKW+VJVPtcUpTQfhYBfiHl2qvSiYcc4+hvr1PSBU6yG
v8eu6jak9iQ636Cj0EgppYmS9LCn7aB/oIfWdlxPFevHBXj1RE76SqO3zYzjRnjl
tSAauTb1pTsxPFw5HJ45/5OwocQJ6HWLIkwgPUzsQnLCUg44Hd02yMUpwSIWwe5p
bjrS42jrB7wwh5kNiW/i68/kzEOPBDhmWjecDlO2+gX/Jnzq3hSFgx5C7g3ofR7p
1oBOkGfD6nVjF70BeMCzuZFWZBXAcRlVS6f5VL0nOUVcuWIc5nJ9Mdd/qpAYwMlv
Dx723frjII1isRvAd107oM7+4jPJUu94134ajxA7ILieuRhnVTxk2rDc3qs7Tj2e
Z4fZw4VmFTxKfmpyABDfSNV4EH7aB4eS6I/ei1abjt0t73ne/gxZieaUMdOJ2Wqj
129x7OMlG7AX0KDkWvehY7BHrB4okcxJYOaTft7CYr/ob/VW/3BAEdQJmkIIg/bF
kT1KllkkdE8ep6oYoGcn+gBqsqcap+sBuqO96YTB5SJdWODe+H+K+UX8x1Ui1HeC
QKKJiiwzph4CuKBumaFqSYJlmMxDrUz16pyldnXxiX0ilfGwjqRBUzacbyo8Lpql
Ylq3MwGjSaW1rjAddg9TGPk3nrzz2zK8hzxVv08KjgGfptE+C83LeuvB3pgyXH8t
r3E2L3jVMmcQb6TPHyXvZPiBomK7hsxdAIt5oWp9OMkcvnA32wi5yfPUb/ByntG1
scr9YrVq2geRb/MRdSwQxTpxMrcsaum/MVyaumTnwp5NCTx3PHleGzY+j5hN3oMc
xD8Tje7mpkrfQf4FSIALzSFwlHFYvz/Mt7XIdjV5r5ATGqdJ63UwH5L1WmPOFWkE
RLYcM/Kvu8L3WIGy0C9dJfWs9RaQ9V9+3UkDPX5APJiiDtQ247xw6DlKCS/RjxfT
GAhF9jxMWANIKuZV3CEc0NLEz0GFhzNOOfsP+MEKPUEmrbDoahtcuLkUgGi3+EJY
m0+U3IDbMc3f9Uk0x47XOc0lDpHIr2UIz7rLsaS2fkOp50s2OblJUeC7Bz4I9Yh9
ZgGbrA2q8olhswpJTeHGpS2WbQvA0UKAcJjFzXIDhN4Cmm6ezGG/Mttw+Rd8le+X
BZdVALbfRWR/llKQTUBwTJZ8rxec6+bOlhOAOICNekW1fLYWL1fjvIHTEFcPl1t8
ffLACAt36SYMeIQuE+V4TCyW+/dINFyXgXubAEcgewCk7Sxs5qb2gNe62PJaokMD
aI/aPfWEVxvio/8r2klX4aJwT0UaZs6P2oVth07wEsl1wKlPxcXJQ4vQyV2ZfrbL
rd/99iArS7aH/iVz0Ykjwbdhgd69QD0i8/Oj9X1dmWHhBZ4l5wTb/wFzhyGLFvf0
P4R0ACn+xV1i3+Z4VJHpTgaV4Weew9lv+8Mvfgl+kSj2R+XA1/bsSvweZ0IeZs2B
5gDWQnFrwjCYqOi6VpTjVJ4fZx4NNoZWmuM1bon9BWDui2w8DxInDGSL1M8PRQnw
ehznzq51963dfGjjDFaUFL1OY3sMLOBI6DE2WIlmpYqig6ktsJl/E6FusCHbYxkl
24ARL0bFDrkARn0PGzIe+aR+HUV9+km70uJhP7s/Q2PBDlQr73jJgfaEtXR07MFz
qa0IR3wiSLqwSFke1yDph0NqDtPl0myTjBSSc7i7wJMjBuw636cVMIYxsPPSZwav
B76Zz6Tgoec4+kvs2NrQ3jZv+KsyaV9XXL9Zzur4hRLWDLDg07OWjGeye1JC6+4j
mSAUTj5zGg5aZDcix/8KMdabXYNrd+4wno1wmNbAG4mvK4DWbcWwHiKxubGbSoc+
bne2udzTJaGBuSiPi2CIMiFviKJ1U7sbohxyOdi2wjQYjPmdyz78SSFN11SyJlYk
J75+n2xu8dgS4moUqahoSZdYWoTvz0WqVHd9AAze6MmohHB802238YK6nS04TAzl
NGlPahwwNa7+/zfaylE1OZqe2jQ4/IWPCDa9hGwwhtGaFlWFNxJ84KbzJkTHWpyc
cD7ysVBBpwK4ULjSSCyBh7DwiUlPa80CxaowTSYZAVudxKrRVBJfGaS+NdJsqPIb
tTg3A23q3CLuDQJ7/FOYMVXL55huRA9XS/2vIzwhJo7GfNGW7OLQOonWKE3Efra7
p5PkDuGxNo0Kbk1lqlhZ+KVqc3HuST7IDggk3n6/1wzUfUY4I1W4vJsCTIUG62MU
4cWvDpCUQvovQWLPL0TocOmvhk6kzsE95N5JODvdztOdftHbVRbaDenix4BcsVck
SZ9dzfD34UTQs7qfSM4p0DtJJsq3ja0jRfr9YShpGuKe6jIV6Rzj5LNa2kHbSYqT
Wad7vAPs65TOt5GNm//NFhnM4kBc3z239iP7Hr0VGxZ/NoK4/D2iu/qVK1mgOAyd
WXHTjAgm6RFAR1Io4VisSSVox39OK+qecT3ZwbZ45l9NiIlureA+VyfkgexVkDa+
+Lep0Do33RtwRTHS9/N4O4hl0mx/IQVhNlT/9jwweQVgGZwrZcfQMRpEx+AFOZBm
9l1tFEIZd+FRZZDiE01r9Pdn3bXur4xgBxl4hok73zZPW3Mb71fcjZWKA0V+RS3U
vrSBtjnzIRapwzdiJhdZgLMPbIFAHU88cqK01/Zk5Gf6DfLmAfg6koPPhMGPVnne
kLrUp/giQkewDqFWGPhZWNSzdWDXTRWQaMqkDWeD2Pp6391OCF4BIToIMPxyYTCE
VRfhIh8i0sZ6QR9xQqrB0CCVOGT7RA3C/GxUzwJQk2AWVsnTEzRmvirvs1hKD+b1
VVxGTBTfjj8DHvAwHbHgs//DIMI4V6zhQG0IrR8T54bYpQ2YwhKcnIbXnIqiTP4l
djQShFZKaUO9lZ1nhv4GIVzS2uModPE7bSSWgRiiJFWXaaI1tXza7jGV+5+epXY0
2X7PaLB5n1K1K4rugOvSyK5nRT1cLzDzyd/xUduoBAeS/O2gNiPyXUuTzxUUDXHp
QM49pYsbcHpNOGMx+Gsbli4/1JR8jh1hngT4S815sbx7qwR8h2NKjTtAReRlBApF
QyYKRp+g77AFp8orwlRkfwgxgrXhHruYVjUmeigKPxLok+oTF5OFQkktm0xI0F8h
jPIJiEer9E7wWtmzKYvZneVy9L1t63ty7/1xDXgwUYeRFyRifCsKtlfHZIgDSLgj
77Tb66qg3HGX6RgW47WkQqPs6SDD9HBigofKfda4FapuIHZKiP8BLfiKKB3ne/1c
QJzU3oNGG7TTb1IaF4ID/mAoAQgsm6N6lE6k4YLOAMXz3h44d+jqXLcL+yp13opT
LZ1tKYMWTyLypvgVCtAbE+aqxvQlmrCLmiiNblUEgjUnXqZX8HcouXBTjsiFEmMt
YNEtifb4efMSgv43x/tpdioK87ub7O/ZmHckZfmJkrlLBnrErqXLiB4VLgJ8dQ1N
wLRi2ienzT8VW0szzJJ+j5NzYlWkWHHU5gSYt49WUwLi0RcrO3I7HZUSN3SdTwkB
GTP+zSiSiKYe3B7+x/5gi+w1qYSVcMXZjGXwWSyCEpr5R5DqefDtbc807VIteK9s
++zbx7BIVdvRwP4W9n2/JAJ0BEmusQUrAhCv1F+ZsstiLWprT/VpWAiTzN5/6e/g
7CHEyKRoTISxfD5s/YdGEm3TdMBKKYhyPRDGGddwnXCh703xFQqKZkQ3EXBtu4M/
PBb5efhMLdkggyEN7okRiSc7huiyXSOTAsAE152PlTneVzThefYD9HXP9+qROYPU
po8GpqKIJcnjTUHJPCQVHt37scBw5uSPsGg5jYU4hyo7nJwSaVyJ0AUo2D4cY/fV
ML1u+x4xzy6aVxegEMbq9tdC6oYwsC0r9kmpPnNUpB9qvPA63u/03yOm6GwBlG5P
PJAuKHWQ09+H0eK2KVWRaUB3FF2cYxhn+4IGjCgy/710VhV4Fx/zzyrvKSStXyLu
62lcrwXZ9qScJ05Pdg3fTdJ58CCkk2zxelxz8HcHG3IWEvt5iz20qXaPOKO16W2+
qbtOAPRqB6lTTo8zYLTNnxNITY/MWLjKy4hZlldlbFM+79ljX+54JByG+W+Ospz1
9Z3TKZ7Zj9FmsydV+Vew7HyUAM/ka97U4+bHRDPAACl0wLQlevY1G0uL28AsKIo1
JD2MpnxlMAEZZ/f96hgA0GY2EXE2kwreZsueHqlmvnv5O7lLq56aeP26l9ijeIDr
lgxILVtXItbUziXCK26dZTB3XoMGmXYg+pzo7u5NyCCSapo1voXFdMF9hWXq6bKo
C2/Vdj4e0FIxbTjm9U7bsE3950AUPyLExjwIttIYPKEnGIoOlFpzLzXqUv2wWefu
dJ7rdUsZDBhIkGA2vw5joQQ/FkD+0XS/xt3mrnfE2K2g/mndcT18puN6g+pZMLbi
/m0+Xf1mHpL2CJf6RSYwJ4tBwflK81LczFUBk4o+d79bI3QsNNzTMnI+lQq4AL9w
9yK5yB+iy2RzeB5H4/8pl3pgjUTxvNbWZmV6WM5OtqFUdcrtf5cEmeDjYEsb21tu
SpQsKOtN7KGU4TB1NxC+EIZu8hznzOJf4/orzK1SuWFZf+4C7gTn85HAxtMzH2HN
0W5VCHQqLOnW0+udgHOdnzmEZqSwAqFHkxdXrgS0BGo2ajk+qIO+KmaFr4dFWjt1
7zbNWHMhwXG8PK0qC2eV8gWpc1kMpmugv4VdvC6cVeNLaFQPO4ug0yqd9ngBtgzW
9nsMyqlpozOBkes9ws260bgVepqngvJ3qy22AM+R0VRCkgDdJcb3+xI/Act7crpO
fA0CFMBHiAyDyWncLLaCf3L2FEKcoAu2NZkAcaRqR06fb4L0ijLK1Zmn64GGtA/U
28wXfe7KJjPlMj+AoH3Ki+Ou7VWPL41WESTN8HPBPtGsQZv5gzqIeVN3hSAUT4QE
isfgEplp1MeqF+cz2ZD8dAk9POeah6ZBIwXVgBAH7mx1JM9RWOdr77o1B1Jo3OrW
jXGV9KEIIo238+cbsSn9Qg+AT2oT8yrffAVKkn8bBkKJO5PTOaFfRaZ2RK1muUet
XmNk6w5oHLjwH0MAo6ahv/hqOtg7N/6TppHUxCvt8oODi5aTCNBPEv4D+2wJ0xJK
KhgSo4wPEuFZ25L9sBvbSRS63muICpTOljfiYGro3yYyY1wFtRQFMEUKi2hQAiYq
8oDHEK6GFH6EkAWDA+05UJ7ZGeTc3kpG9/TlT5aNLsy23oikPnpablxyd5j84OU2
2LiRsWic/pXyJiBX6FNLr20dTZcobAkESNabSFLF5b3EQykTVJqetELeDi2Uyjuy
7P05oVoM9zKDEEhZ4QO9QIpfBZ505Nktz85eF46W5NlUXA/15c3PA19dbiAw3qE8
gfw7o//csm3ropjcqrIqTqI/ia845jtRRyb1tr2BWNQa5UV2ztpVB19/5VHwaLel
gNbE7CC1tqRYyg3JTViIkWnq/Uhizs4SqMkXu5m8+/n+Y42VbwR1t3dDaNqC6VEV
IBYdFoyd+rZTFGSJI53YtcXXvR9/8k0CM6P3+qucLKXu7L4EM7MWDVrEBPKiF+Ch
eq7dnK5Vudl/qlAyxjx3YJEQDPsTSlXPBBzh/XbLkS8AydyNsYL/Z8LpQjOcct3/
Ksk2L5SpXHBEB0HWxWV/2GobzHmlf9PZOQ9vHbQlBANA6xgs27AHBDKzHYcsm9EO
1mHjtF5izIE8wmH6n3V664Xi4Ylp3pOq8Pfm4nXBfYWizL6VG3BmsOnI0xDCFZtg
eIl8D/BSVeo4vXZ4oowHo28XYvAaARdHbzWnyfeJKaAMG2sHZwyL4VLDoyJBUGK6
jsuMauf1yDAT6Srfxl3qpY3VdkRcgfK7z5gobhwyLTUARPOZklEML1Cpre6sL6cq
KBODn4wMNbd53tHPz6L7hxT/PMDzYbXC5DuWct9qY1Bnk2AcNz4a5z9YrD2iX3Hm
OkVdWBqobxQix3d3RwyLGg33J+X/UNl9J1DGZMAocy01GAYEXnr7bEs61IkVFAxp
4FsGrW5Y1AGm60+ZxfPcE+r3d7OsHEbY8O4KhgXB796Y1fcwudaboc7IcLdjoaGz
ojUPE2aDd0VvmSieT8w6a9h1UYKZ+8AgWKkHln5ef/lzgh1XW+ZVMqjWrMSYHlJN
76mFiSd3XRn7NxoQ1Ar65FNpIioh84uD1eSNQyLHCFzSbARdt6HtUicJvD4Ef0VM
q1HLdzACh9h37DiJLTcdnXuXH7c6E1jwQXQnTOChKf2QFZT7sGQuA1HIDWFfu9Br
TknaRjdru5wPuzaKv4hu55nTBLm+ra+gmIP92QicOBh8qPlmONooTYpl+EGvM2dU
gBMdr4tWQy4LJs90vB9owApEbu/3CTqVnAfknZkFGV3PVgCjJZMmlvzlrpLgJy76
gSlcGUVqbppTNQVW0rXEmgXlLp9lHC3kvg2DzZ+jCXhLCRV6YY3bfTo4l/TtFheE
uHW3FQWUHJkhC8FAIIC9oOUUbGv6eynR4gTftehR5/cf4s+pwCGG4eeROmGu7Lm/
7WSJJx1qOQb4MgdKEGvQsO2u36cw5d88WzDWPabMVZJFOjfSdCsGAaFcUTHAMqJ6
+3d/A6m2rJh4J5Rh4Dz8F5OWqEzrMjYx/SGxCluId8LW/5dEMexWYPRhIExIlza9
XAy36PzqCoxE8eT0lCdSW5+Hl01U99jHl2YOs1tCt+C4EmkXL6lnKZnwuhbOWDcG
g1JIuwLr63oGm/SzfK7z3sOz/Zq6GXyhi+XvdSwYa/wxYMDle0kUwr12XEBmXhXJ
4lP7p6us37KY+2jR1sd1YiyiwvjtkglPxLfblv9HUyH1tb2IIXGOkyoCirNsuVLv
r5SWWfBIoolh6VGkEvY+A3FDBmFWe5K+8fORFri1Pj9PIWfTbSWJ95AyuYNsxrO7
86Rz6hZgNpasOcB13uHXv2jHrKNvOAEzS+J9otywJqjiD1LyiQ1Qch7pj8VJt7i1
eNn+D0HG9SC+BTc02vn9DnQaHJ9C0cugTIz93Gn8jlUrXYuRAAZ8wtS3nBaaU9rR
A20Y5k8AdtoplWzI+cVJ/fQjKdXFHaV2wuJxFH8v44Trduca8AkO7YmneCWEh5NX
g42vgEiz4ShKw5dqKa5QFcmDtMVEpYRK45j6GYse7XmdXEOxyS7YP7HpkKH8xSIw
qaZIQH8S8hKrqvNCWZJcEGnlUN+21Zi9exG/Wvfa0SJSbuFSb0sklleVQCG+ot3v
8xKPc/su092JH2wcSYK/QXtWH3WL6j8PXUHsubPMi0sit8CXQK6Bqh1lpOzXp2yj
2/PRclA9zAtXVlkGPpav7h9df6kqmPl6jwZt5Kxq7inwzFAhT43DZowEc5zuJNzk
+reBVyWaN1Dg5Dy9u7MxbVAijfsLfHq2EkQspoYyxW171XGWxJTGCn+hGUI4VlsG
Zw03ibbKZrEi9B42BkBLsYiX98dIYLTK6395rTZnNp8+9ywYOdGK0uHqO3An+QJn
ZrmUVQ8mIemYQLr2Skp9DVm+oHeEtCsvpFXj1xxuyQmuNv8bG9/QYh6ohygV90SU
n8cFa1TDV3Nw2o9smfrKL6as6R18/TwHNVk7vH4/F/L9L+gfL8OCAF99YIA2CBrQ
nst5CLp0wLzTT+WSCBvGAF5TXGxZJeFSTEpMCGx9eUpPulesgwS2RO6zeGzKPwKa
VGPRlIOjkRrkMSnLMtWkD0fBNkcfCAfHEuk3VbApE5mHdHDjjOKirw2TolB1/qQw
GzajTpx0VEPON3/VF1QRZ73kDnQR3kdaPcK4I2To/7E4SzqvPKZSIW1Mt0PsaYi3
8iWxwSklK0f2VmLKN863j2N6En5m4L6n6l2xGE6DW57AgqDsrPYUn+58+AHBoNsV
5FrxFlDZI3vxQWh+H8JoMnhK6eqG0ZeFOCI2RLip20TzaAhNt6S/s5FAM0b+PYuM
HsrFmlF6Ih/ywR3uw/Tctm0kx3Cd2KM7attgI9BtTVtnz9DDFgg7XFVwk+celt1e
oxs5bBDCAUuOzkRRG3APbU1eBbZ/joQuqsDwNJcCF+MGy6Hv1UwooBdX9PkjgklD
AjmSkJjVneA5PS7okN0oSCRDl4lLsvyPPrc3SgWrfrZRlTNmIafLBpqKo4zrH46S
cUKmgCAr1O9UCcVz5FFfcQ9QiJxe9xxVOhDnIqGAoeUXq6Lpwqwz+R/IcPVGGfBL
FheUaUWwDuIc9x7e8+FLl9XcSszXWCePcpcFlpiuqqKP639llHfvHzKFprwUGBNO
zhYwf89UyNoB+lR+c0bVL9mj3C0/Xxkv6oQwAQiJnkE6PHYJkOOc1Kb091uLd8+W
AXHl15abktbLQohZmDJ9W0qqSERa3JqmC/2Zx2psQ/e3vA1FEabwvalogt2FeJRf
GzBqqHOuCZFpIm4/skvHo7JlggZqdA6XbRhuD0ku5t7MAk1ZoOu55f8YswlwMKc5
2Ey98d+Se7aDUQpu74j9esGDjBlh0x/8R4XG1jp7xxDZ6sjgTNcYEgv2ekbDps1p
zwAKYwbm6PEYCNKg9pEhnXXi7dCb23VvSYXHQIPuDtzptmiqRxjWT4efm0GVQkgC
jAThANylRPLT3xwTYT42kXF9Jo2XcuxaVGgNwTba2CN6+u02Bw/NL29oue0hAJw5
/x1/NOt4fAO/63FTGXjGhKEIYggiIUIIfKA+bIn7uvEUVH0KgaseksikGDe+W3QR
/StOXNpUBpIHt1sZ74xXqUpHB4jKNKz+Je4C/aVUjtDrqQaoVYrNxY1UZaBOZsWg
xjk0T90+V8vo+0oiYt0+dwO0byeQJu8rCVf88hJntxnR07eRcx30XDaJ75Bg8eES
ruP/GjitmgDCdg0XVFhususkBTQDuvuX7C/KNJOVEpktspbwyLSv8c7uQjg00Zjv
HqVHLfSZ6drRb+Y6a/lrm6SDt9Idlxvf8Q+8MA6eu5TGYvre6YcUXjPCP2FQnJLE
rVQ34sDcyxQEiT6+X0sAN169vqqVX8fM31wVqYJnXmvHivYRlolSR2i/maFF/5EZ
NQi6du6jv5IMuAkcyShRBh1t9hz8x7KcWJvmoxL5u/+PMACSQKyU/f0tnu94CZgI
3BkJ8iW8kcw3XFjJIojbJYC1CcejSrOzN1Rz8tkqKZVjLIE2uNx1XxJWbjL8/lS9
ZwCujkwUzoQuRUgZFb5qj3PFJJrUNGbEoeoKECi0TKHu4X3HTa74y+mQ6dEodrZJ
UHsKqCa0YPTj4FM5549EYHH0O/0cHgGyZFYGlfdWVmkXbGgC3pZWrwjPbRwFw0/4
9n/K9IKcQSAOli+d+5X+b5K6EDD48Q0+LTerkbvECIa9EH7iNaGJRftxhudPvmoc
Tsbw+2ehZubCZd7f4yJPfOadTCcUGZfOzfYK1YxxDDtS7LAXFO1TwEInxN5h1SIt
P3EQAv3ZbNhCHXrUOuX62oAV0fFxScW15LNfscl08wjEg0+KwcY5qyKfOYomnGsg
JoYmonj9NKwVMJDiA/BzrhJdlEVVPqfn3zc5XvHe2LVZ2uApuN6P7eGxqCmuvUwg
j1j4d6xjU5qLtKYej5cxqK/E4/ktS4LjVzNmskv/8H3fefP3BCsG6kAspAiS5RXo
CCAlSv7mGyYSZ1tzk49Qq0k7z3B2xd62OpK/hXr681+UwfDn/s8mxcqvo4ULMvyM
NbULj9I2fRgbbpYpaksgFrO3j+oZudTDpVXE8wLsaKHECqEintrd5tx3fn8OKeQU
QCPZXl+0oOH2uezhw90yi3RMuB2wnTcYUgzfIW5Ntx7Qw/bS/bu2Jzpx7ObAlb/a
KxAiIhrlQu+uWAoFzumYR2MbIW+l6aXLVx6TJyzE7WpgldeysqhS7B85UQm9NX+7
Gt1h4952mvjMUGHxGpg9Ia6c6eOnxFQB+pYQvZJmIZ9M79OVhnVNj2cUyN2gVoqB
VMjWz3C/176V8Be+AM4xQUOHsApk7ACrybLX990OG3Fl4/BroudI/epsgk5akLVV
HPmB7OQ2MFUnnsnAe7v9WipNGMVskYlv9JV37XICDvDKQa4ots0KxjeMO4wT4t5/
dvpjmsZ6thWeTMjfRDAF/JF+6YunkImohQXOQ93psFgXvcNAdMECChIztYTpsGoo
u7tGiIwWMVAeg1nUmF89V6TE/lddu5kOB6TqvHUYQ6GhqMKxkfxqrV0BOocJme3M
+EQIBsM0l/JtMxG2DmFitUkVcH0opCK7jNNtkm6x2AUdssDhd59IF6bggD9RBGOY
XuHirFQtbtGbTeRCOqBoYWIenrN2SdiDzJcQ+gXncERkiJBgPduymR0hXLroBaKp
jpRKRFsIOpT1wrg4ffxErc1F3nXOtOORMqBNsXrX/Bb6Bfrr3HFKuP1jC81DWaEN
F/aFkMXDSREcSp3F9hO/J7MfNUV7je0PHo2l5BPGNJIjw/TVhLDIl2JxgwttPsTp
1W01yt7LJeBI7u26ccyx0ul5CNIB/av8P6cll6aBialLBExA/c5OI0mRQGTAr2B5
Z+RPyexjwM8p1eQeGhBgV0esG0shYbm+MmJqT1Z9lv1JKHCNYNAAhyrDNrQKjRof
/0tdaMDL78C2YfF0Hj8R5otCZkMgGZYKd/1AwNeISgsDWoji40jzyXaI+Wl3h0o2
XMw7g+mO+WZaUROiYdn5uIKvkMvMmyCB1IuLSC+bEL5z016WsvoloxkSMda1fqyH
7I8VUXICSpcjUQUjs5Pm+N5bJn8TTteXPh0ByInEGmaVG1FUE4Jv2GRRByQFogsN
fp6jR5P+GOv/lPfwK0zzTu0jRjwqWHUqD1iPE/RJNNpjYeEz4WUdLpskiKd+RyGw
RvDnzshEyzyC2inHhiTiqVf94/ryYORBKsVrU+V8UaAMmjq9Ha+LSTzs340k2T9y
cEcnCeUhbW3BrtFZMlOFu0cUooKtpGNqIfB99jr5r3ppaG1DqPQr3whPlw+y5T1i
9rU4wCuce+LC2r+CEzsDl0YZ2oJOQIlCph/tAlzpLBSofYKFSKv3NdyehHrpuwo2
mgaIIBAmswWj83CEUkhb1Qi6zFnHdEEngw7RZv7oU1rnlmJzoQhICv12+b151cgD
mrbQj5KIcFDHdco1cyiV8TLv2nAoSIhfDmF2ZLZ2Sr791Zevw4yMK51Ha+qDbPVM
V8tsuhygLbOSXeIPIrGD4SNJ3SjWpMZkqsolAXvgZ6DF02kbTyGHdScOy3XOXavS
puIxSfO01y0gLWwifhzcMwxRdLNYlUFYRaE++6JrMuuHamw/StUszQPrcbngYiWh
kaL97P5IATxu3Ry2EvThr5jqVq7TcHLTtxaHaOwYpSr98pjzNx6Qcm2S/zqDCj8n
5oyiWa1TzdqEy+8CFQjvf16MXSviIp4H3dYGKBHLYpw+OvCe5fqUf8pHsbYvCLjc
p/gGZ1kye+a8Wv/j+QHPoRH5pTSZgzUyCTXrrROQQM8+woTo4ZefTuGPIVPmWhi+
rUsRB5ow47XJBFBaSErsOnWL5hEO/XNoW1u2ptfBsgxbEypsKBa0daz/k47AnhQC
ILYsX1A8iY6aIMCnseLoTzPx8208OJhuTJIZga6DqlQitzgRuqpKv3iVuO9ZfNNG
UrogR38Giqzz2PxC7F434YWDPoGFeHyLq5w5A/V2Fap3/ltNpRq/UIF/IxhrHlWx
krroiM++RES6e5WXiT25L2CFiUtipE5xcT0/FF/wtyzBL+Jb3LKx4L2Wszf6YePP
VZzSS5Dj/a5own41RN1HtTY5Xqu+8zVHuzPQKtNeVHovi7OmAGKsJdznGmsa9tYN
4ChjfWgYycUfJy9RoC9p80NrKJDzfa+4xCXGiQDszixG3oN6jX5D+viIxQs6zftm
C+4jq1wYEo4/bqbsr+YA68jlBKf8kuuJars9QohsnmuyLoRVb33z0KyWwuefUdaZ
6aoY1/7AZpXwCezLMPHDGa3o16+/2uHKFcYXQz9NxfnZcIBhRjwn5aWo4gbpnmeN
c4iJjTEiMXX9GDj8QbMCTATCMcr+Yb+5iTeGm7wu2e2MtvE/SmkLG7ML0NA7U2/3
oPaWYbLKaaLQ9g9viqoM5MrrQEBJ3AFHekqo8oeyCfcK1zxbzWN/UoEqrFsHPBtO
5pGZ25LiW8inxqkjGXbgpWv6bWngHsz3goq3pCx2lafY/qR47jC2m4XRho7jd4BF
v1Y1M8s6VimVXGTqpIc43FDb84s1vcLtQHXFTJLpH3U2D3KwaLPOBEvrPY/+wtYS
WTfOZ6zgATF4ezsHj4XyInLhrF6I1+YG/VMsAxSXDhSF4XG4Qy228aL67WpPnABO
81eTl4zNHar9Ui09Y+9QQu6W1N63KpdqZ3zA1xr9ZUYRReNFMn4hUe2Fk440mB10
tOKgmkt+WQkGoiSPld3DgIgaR8K42ZUv1cSMhRwcGcOI0LC7Gi3aI3F4TE/RvH1X
9dmJ/z8W3jEE5TLM7xx80p98cGVsHCOdbdG4aCRdJ4Uhiiqp6+7JezFzSTDHt+Pk
tq16WCB5D1WC1IuvTV1hxXovQGvrmqBSw5V+m7oyt63Iw2cWlZMwt2kFQuxxUxwb
KITwJnO/wICjUdk09ManyPfOjhgTUvxU26jGFYGt8uyBY57eOeq8HUPlzc+z5hQ3
jpEQ1ZajVBcYGdjJvlJqyTEk+rwlto2iOH5HGLFV9TfzoezBmUvk0OxMp0HggwqS
fld3XdVOblV3FII4TLtNFErTJD/iLyfgIv4Iix3WUcH7pUf7aknbWOEYclA840kK
GpsaYahol0S2h6JMkdH2Kk//ie6fO2WqS04TmVne+619Qz26alV9AiCLBGml7uVN
ejRetjq1SelhtiMhxzlYPj0CmRYjzzGMdX8yKEhJt2ywZ74v/2ZizuGBneZh9vMY
Fce09QsFVjh/Ps2lhFCV7Y00Tz9XW5EyB7FmP5iEN+RS9158sNRG31HaHVDXRWUv
WxlO7iS7tFTlek9M+BAQLonEuD+Fy5U3kvl8v3FgvsQf40lpqygRo5xg4Jg4/UGN
DOTJcqecNCpJfdC3nLYns0apJvC2LABZg78kA7/Z0nbny2UxSgxSJeK4giODKdHH
YK/MrMg8u+cSYwvYNculfjQFqMO/nkmLWZ9eA3rpc2laAhHNhKb5ybIFwu79HbQK
2SpYV1Pnb7Azbpkgqkl3GjNgDu39sAYmdMEnESs1eBzQOECTTydGcWGfq8EoCZ07
yEYeyiVna0FnpLdGEhKCCFGh+wXUKv9JmktqsKtD5qJsYlQHuKW7NbTwyjrGqaCz
VohxirxSAwJUuhCbcqwKPYgHRvgY0yXHsvImTK/wVJa4i9gGqOrG8pg1A6L+eKPh
Ol4qWZy7lTM7KEATMq4TuXBKSBn+biTgGsOBSyQoekJS2zmzJnnRj7LgHjEceFE0
wFLKlLjgJu5Qzi1MsBrUIl+UFLySz1SbSiQQcVWMFOIyF2JMxAwuXOCfqY2qtWow
NPkPx5eXkTannr82VkSNNZGMqmtnmrPbg57FyCKZl6dTASycQ7CGQR1xTCteRl5T
gGgmksr6j5qc8DyxGLsDl6GKQLy2SAx1azINMDTnzGJOU6jvkRML0Nj2Um7BTSSj
aumtkivfJgnM1to0sD3XWQmRa8IQzjFgbyC7xzn5ky50iubvhi3JB6oIGrf8rH8Q
8TB8V8hIbGFaSnZVsHxCrUXO3ceFVXKBshKUDaQzl9w73JHK/pkgwUFDUrB9gsmv
Vri0aIryjBnxPoioHSqhaI4oJ/HQJRM10aSf5fJdQyyWiuhtmfIG07Emcbto+pEm
HnHrrxCDmCS6CYeR3KM8KAcO7ZuJE31SjNp23+SjxiUSCkRr3eyVSI3ZlnCwU2Ot
cNYlgaMC8jvRzjOKIFnctaLUTXsz2aeOMjlM64OXjwongSvFgj/78Bp8ISnN4jON
bRNV1dgfwGg0/f1t+4+5Dqgf8zwG3exx7KK190Tq5lNEOHWzLCCamqokQ5ap2MTl
r8l05nflzfqpFG60kQENO1tVerLcd6nRIFY+1aGznrhfam7C5tvvIFVX6UviegTu
+pdwry22TNB/ByCzQP1+lUwCBE5mw55+78GbHyK2iJhU+VaLRzloHbMG8LRxen7E
BZbq5/aVoXkqbuhsVNHvaX7kabkk0EHAgpbGmduYkDIzwcmJ3ZswdYJsW4fTZiMu
lIxmCzOpeloUVSgzx/PFYCsljdXWM00Z7OZxyWMX64wU5cABEnQmtvHOeC3Fy2mX
QkDkOI8tP+DOIaCKMFsdTTtbLrNy7PRmb8bjuUtJcWu4NQRQ5KrqGfXlQZhvoB66
tYrWq9aew+jYt0ty+rke5QFfqXAWs3yJjcVkGTpE0DVzlGJx2ROjTRTEeneZdpS5
T3Y3zvaqeUrXbbsELfyamjKtz9cs1xsr8ER9XEYpGaT8zanOzpEqQODwIKFs4s0g
pDhDeKpcnJ0W9AOXSAwNHS1736cRvOyTfzUSJ1KK8S6sOJWzv2SlQekZ6QNqubxC
uLrrcC9m1hSvHSWgXBTHeFZWZxu1rF7ClbYWNo4VaJTyf/5mlo9oH6PiEaZG7tQt
AanndJj83txTvxG9pXfORsOdZ/1I3Qck6LEgK/9wIjW5uq1V07BSMZX+1HB54GvT
UfpCufdzuGFzIy0kz7r34pXR8H0fQWq3gwCNZMc7mivIff1MrLGQEHNUbZ1FtMWr
iXYHaBTkoc4HitOdTSNAxiTSkU8+P15kuhyhdt2d8XKY0Gd+Ra2Rbs4SIV8vqja0
cY+iFX0QgwOsCUhP0hH3NPE+oxXh+svD9Vve461eXV5EZhP/1iOhUsflj7SysFs1
DtA/aDnMxlhtrl+D5A81F5/sR293WzttYt1ocz6jyqlvdD4qqGdP1neh3rZVrVQL
QacJnvcFhdf3dv9iSG8HsJ0E8OZU/dUB3X/S55I26UZHRcTXJ8efLZwNOYMHUioE
CcA7yhTcaRey4GhGyX03gcUVWe7TQK4VHqrOL7uns7VgSrvgHKY0OxMzqgu9kQ1F
7kikQuTd72lVeUeceVd4PsFzs7/9nwv0THPV4eWMdKyROs84nu2JUuijIaWnpRef
QWmX6TlLTQGUbHwZvIChRUXL0OXYEeTPRhcn81h+mB0G6/gTWELtY+RONsxAgVXn
ZrSyzxPa1cS6iCaPVKjwNDk3FXC6/SsCYKh5OrkyWPCFKWbwOU08wTe57lPYSqsL
iexF6j5L/GtitvuE79blmPwO1VxXqZCdilYSAcHglfBizils+DeYfOsOLaH8kfXF
LHU3riyvflt55+nm+FRXOfaIJfIKvNcopQGiFSU5cwBi6lu3I85b+cU91lYrjs0f
WqWVtrijWfN+PWlVJTcd1pm//vsHOZB3CzsGkjk2rWlFLNrvN0DyVjdazLxAhlY+
WdNQaf08aDKguVKsaXdX5/pnQS41SHNxCAl24IFYmf6dSl55zsJALesI1Bw4SuSV
PJLpVl7WQN7sRGVA9ruxR5xIvgBDOehp0D5uRu3ud/ZZs1N/9xCEsaglgr6GCuO7
T4b+ZJ2LDsFRHgoswvH2p8in3fOy+Q5vSpobT8352zCOQi6TZprw1c3yUxlSxWOH
3DfTIpVocKebmjU7KPreaaFZtvkcVvMT31HJMwC2uPLePhowBHR7yZq71ODxxGqf
FM2QKZlXpESkUWK1oPxKulUREBs4XS76zBX9MPhYSJa1BfsEcOUCa3U1L+fD2E/f
TJkS5V8p5AD1lm5JFujbH7ZD/oekYRHYVPs1GsA3c6jKADjtLvhDJweHKPvuKYCT
WuScfgnzf9Wdl/7Iz2me620GJrqAPme9j8q/h8oBDlZ9eXu+wNJxOLw1LxMRcvns
q7QDT7t21MaWtZNWgDXWQok691RFWDDd/yOx2yMIhUFMKm1NAqmn+TcHhGlLxth/
R9rzEKFmuKNgw5nrpfwIYRS5dzErKyxRkS90Q5amC2RblLYz4+REcZE3ORkQ6yJc
cnYPWay0RmhAJGyIPh3os//kNmE+u5oySEgkjf7BdwwBjNQ19DACKOGV+iztg3Hb
dKI0j3PBv0eb8OHXiMGc0tdL4Suj6ArDpi5pmVuQTnrpsVy3QWz2qjIsKJBJVZmW
7JA7FmYfhqekjsmhPzDDIZf1EHd3vFWpS89HSpCLunSsIce/IkDJX2RVnYcJfWks
Zsl6tYI34aP4d9MOrY1DKn7gsD9zk31R6PDWHsWYaK/ttvEmdg9VpU8h09oB2pL1
9rT/072Qc/xyyQIjNM5WCOQh5MNB2sbXuw0N+0qH3Xi3qFpDFBQzd+4u9obHwV3R
HWYk7V+BdAIakM1m1QdBy9Hp4i5VkFnoC960aP7+9PD8OwdjacoOk899N705rtLX
+G8mQyX0DiMkDUur1UbmgpyEq3iqhKCMIy12TNc2QP31g9srR+o/8VMBMBdtzH8R
DLCkTk6V6rt1sh6ngQCIllqQc2sv677oZf4U1KlFMbi9Kf6L1ETDgc8NREQ7heCw
U/aRbOtL5lMW2/ydIeurouttIUuRzZIFk2vrnFrlvrvQ/rir7B3/hT9VGF/oLU6Y
rQnmyzi32CoET3sau/hFMQOefRx70TIZvcEkORhul7G/P7Y74PmMSwUm3cRA8HJA
olS8v8i39wvEtEw5M0GBa6Qn1TsTvY+w691QQ/t3FOB1jSYUh9lw3UPzoKOe8HJl
WoXfxCe4ON1RkYTQ9t6RMw+PmLgf/EK9B18lbnQEUmo/vFjuO8ri0uamq4mZcy4m
pr4Q3K6yAxCGLpWNavk3Hn/Rh1LFqta+08hir8fwDgdzynYLyXsC4nvDWTDnqQTQ
SwdAtCCIKYzdy/W7qer9MIGYKYoRNW5Ey/juXUI/2pfZMxmo2YGnx0inEu5Z/m9s
DuVkdQybJerS5nXFtdRGClukLe4pPLsNLYs0BS0YVZ/WNgn11YdL8ud4NylYHafV
O8N6wgztR3W+zCCLtq68ePcMtOP+Cf5ZCx1Jhcs9sKC6pMGmO/AzJHUz9xLTWycc
9/Kx59qrN1m7dGmcYaUwTESLO6spbc1WCkMtXztifhdGjF9tjm/z8C6zQoFgj7FI
vYnuMfgYrtoAFVqHuZK0ChRGfgM9Of7UTieLJrSHBIr22xcPN/VS3qRNweFZUUaZ
gvOKZbLGk3DPqNOisQSOlsvFMp6oi9nU9RSHOLt1lqCkUkt15XCfDixFXEpmdltt
eBgs8Yzbz7Oq/mreoO55V5DSvS5R92OJk78ishKGNdlKsKFyr8ff8bTmx+7TqL8b
vXjSOS+tPSW+EBsUtU3NuMRHFtTNt66aFmCUP6BNLPGnGj2yvf4KLv6/n0cKyrqx
ef54FpMLInN1LJWRyGJAajWfbFKq9elsCIK/4Xf485v3PxZeo8/AFzwr8enkN6Uz
HiHXsh/fNbAY8txG/QJoRChf1URMYPAszatxx+UCM78qd8fzZ0pmg9gNMRhe9krD
ADjiEEfFPAXgm0KvpW1CU4ju6ta3aBLBw2NMtkosCWaUd+oSLj2oPGfLK84Y35j9
T9zOrgXcZOo8AecW0IxuumZsp9Jkqgiy4yqqhfsWSIJUQd4tQz2Iv2R0AUHxE/56
NE464G5KFQZEJm9V1XR69NSkmmZWVxYsNQjeo6By3lhG9V+vlSq4Q2BsfggnQi0c
tXtFKo3WCPjuM0nwzGVmOJbghma1Qie0A3xc7y+TMMbCzTIAAycRg+XGOBr7NDbk
VjtYeAiUhhJvflgE1X5iILzq7OYsMzhD8o4gbdcUbUMNF2i4mujOdjDhkln7pOvK
HJdxrP4gERzFRGO/543vVVI+5vlJi1xQgzATqmaHZmkqhjJM6nycRyR34gSqeO9P
litwvc7b77GNFsk+aSZadJu4MYN2HNDTX/V52jmpkHIKSvSY9kL2xN+kNEhetTfS
QsmsY1pOTDAgGbO9kP7QYPs9CL3F5zx8B4whdLtT6rX6oiI9gdtrt7t8sB4M+AWQ
GKs420Nk/TQ0OOKJjCR1zVBZR8UjPexlkMteXi1pzaAJ6LYa0EWmSFc54jSabtom
6iz1OQ/CMKIA+EW8tdchwOA/zUhXReFyFamYvDw4On8wYAyEMieDaqWcVqH71FRl
MkIzXlEu//6dZY40ZHArTrjHW5R2nRqvmC6AiDuqRm4ZJ193uNqnc+jpv/HRduph
jABwmhkhc7jkWhLV0X4AndFXvBjNYA6OZQb/rwHW5rRV9JudRIz2B4cxxBKLiD9V
Sjk9AxkvjwUmLqUq9KjenMg1X37uVVPXI4rOndf1u+VEcauZ+ggR9N8A03HT/62Z
vegzrJ1XMIgo1y4ZixixH1zJyPHNjYije0IIGVFhmrBpYQHkRP79CQ8D5CT7DhAu
+eBfNcf43nP4KZjYbCw2qXwZ9I8ETMnZRcX+tV+PR1lWCJhm6hWMtg7eKM9B4tPY
VJGi08LO0r/O2Lk5qm2vQNk1F2RkMvX2kZ3LRNOK4o9FL1qjqNYMvDax1vOs6MTj
zcXMG1L8XU0kI9ZyeX+9Crtc+J4RZKP5h6rq3XBx+ffKKLvG1ZTR47bpnHMg1O/k
LM4y47sluMpJtIhIZEAXoijaNdVuIbclg5macglUuaXqvl+U2AuzT+6mq0P0oDBA
YTx41Vmfmlj8dIjt2crs3CPpbmkhtpIBQywJTaAzRgTxE6/C1Z9I2idiNRLYgfOW
MDI6exIz2tJ9wZVDufjI5IU/8qLQxi8dmvMMuqElBMd4zrHNhs80W3Z5Coyq6jSx
FXB3OtiGfRqon6+bSAaZdsx3C1IECGkNDGIX13LMuU544MdDUYAp3Y+3CTsflvG8
UFCC9zSd7zlVM2TvdPxU5LnwdXciomt1+/s1RKdlHPwqduuWEexBybg51FRUN4N2
QF1RHFSRoXIjmVWdO4cCXC+PyTfIgk9jFYNvZBMzzy2EECtY3db+L03CbkVDvYiB
xktTNLk+rro1cwzEKpaLl96/q44t4jrzI70oXrBnZ0gsRAG9hWGajAQ5bq/cghnt
VwSgbOa/bz6TWCipNwLdsSbT6XiQvKEsE4t30U3751nisd2RkWk+YqlAHnATobDr
L2hP7P2K/HjDrX0Em6nevKOHi3DSsa9ZG4tJHVSg09x/+KQZc6U+Aw9J1LLkrUUu
wa8cVCt0+eCgP8yLdsujGyE9P+VoYcV6FB0pt4yRkdUiRvKybnEYK97U19onBML/
qE8fBBX5y18Rrv5U0jhevSiF92L/36DQpRn18/XSLLQVgyOvlF3UXo5T9WgzznHa
9SN3yDZoil/Qg4ZgoWs3hUykKQrx4XNNhKv6IV2Fb3B9zjHjS/LRyl5sWMOqI/SD
9g41dWNr5cXOUK/X45Euy9WIcyo12e33oKRUF9gzGx0TeGbojL46tTCddrl5Q9Gu
2sNm8inC0nmFcSpGkgnFaohor+bnPKo8i4Q94DpqIth8xz9HKU4ahc+bbvdNjRv2
JmNFnaJPV72Z9+q8ZEqbh4i8I8xW3jOAj+S39uNWwabGzNqsY5bR9u/VQbT8sH33
jfC/CW98Clf3+w7mqTGfNwUWnwtJvKqgxTpdhT6LA0gu/vpwsZQN7EfW/vNLKbya
rXsUpw+NeyzJVG8KUZ2/PTxcNlNZ8RyutLFUAQ7Xfn9qUKlGYSJ8/awq1LGDPMYO
2mTlkC5HhWZuouScE3cFMc/7FCDlIxWW4/g+twjaLPXX/TaCFMKGJClWSZRYFO2I
jVAIItarkNQpeWVeHJxdDqwi/X3wYNodXJZiYBzoe7jkH/oIYd9z5+X8rj+KLtFE
/vvLPJsNibj7GNZTZT5jBbZTb+Ahe/Jx1dtjHtQ1sNnN03cxBXDedp44UhNbFzJN
Fv07mUMmazuCfhTmt4ryvnoPXqoq/fTMFP/8dm4FATd6Gjz+pPhlK6PXex2yrLeN
7ocezIPfmiZPJeGleACYNRdVyt3iuxorNFIWg9ChOb+RRId6710kpW3Ifg5wYWDB
CgPAnrbix904ozxYiRIr3s63y2sqaYQpashVZ0THliKN8xlnGouhiJbHo1bK4N+r
Vw+8THsoT7vQucO8fKYRan1vEd4clryejXSkFLVqfEqKSn9oOTQs3Pgy+h7zsN51
kfOr96UQyjQwObxgItyCEOCCkdHLd9f4Jd6o3IVaZcylbQcLSt0AiJ70BgG0JOTh
pz8vocrTtpdyNOd1BZkvQGZq5juEBQ/UNPbqACylAgCw54BaNieopVSHXSgdbKKw
0Xcw/jtxUpC9cGPrs5L23E1VyFZnNd9aU/SfAVV5vlCoqK8hyCACw2HTMVW1bmF0
cszd+pnLTUeP9seSYUMEIhPym+XUE0R9rUvX2pGfVcvZ55pApuv5woREp9uTx6Pe
JMGK7jgkCZYWRDGlcgNA5iF7kemvOynkDClF1gcf9wAWwkid2Npc/DclRoMJj89i
NtylMUiAXw7zwWVHi5BJ/kT1de9EdfQMIL87FDBO0x8+M47yGNgcdlM3bT/PwPwN
rtRVc9OQVrtNNStyLpYZLr1Hk8PBEw6c7gozKh2uGSpF1NEkhKAxtf2VdRhfgGLp
vvW+UMrMZKraQpZIY6ynHhCenBZw+n0nblr2Tt7DgxzyWUfEA4NKVm9XWScU/u5v
ufKHhbVPhFNkNwuDru/o2zOftIuXk6auws7ud5df+IWAI6b/pqXECbLW/n2qEo9m
SKrqnIOWMmXzR/GqE0vZ+wE1ZSPcmlw8XvPZRKB5qoIgwWAiduhGF767fG250d9O
yonoWurCulaa4FhxK9X7zp7hYGiuf1yVuQ2hmTVKKlNzAhyrnitBtmfpDFx/OS91
8WLfWYuQuIb9MY16i7kU7vA2Pl6crw7I/XCQ+i7girZPA7jzeirTwW5ugoOyxO0G
pDBgDZkbTWWVSp6RZXLtxZ+b20EyYDICaCsUXToe380K8ZdDvJpYdbwgYJl7hFdJ
QsuZ2zY1Wensf0VvCNJgwulXLDnmqbmcFE1Fn3V0vhts2tYeV0gNhlZbBp+8H9ik
QL7SZ/RDxtqhCelByr0PmZtAIf1RTESdJJcKbnUOezG0iexyit5xZtoE19ejL3op
mNo6Dzf98taCxkN1DN4h4nWExGVAlScAOMzxIolykpGXLu4VsV/T7xguYZA+wiDM
mrTt+2usyjOw2zIFI51AYVhMIlE+ilqw70QJMXkUMvCY2EDcHflHzoUv2BnM9m/L
j6FzlGOjTmZJfB7XKXP9OE0JC1XIY97kLBsjaqwCuJfa7lqdxbC7uNsF9mDtCnxJ
YNio44cPIdFtzGpthM3dS63Da+e3kmQFqhg5jm03wI+ikGYATSTw+dUO791y1GAD
215XC0jW10jvVBbL4r08+dzzIgRSUBRoklbA6gjE8qLvUBc3QF2yQbytYJihx3AU
syxcx8hDP/zAIKhrOpt2fl5z+5oTZt3ZCw3MpVmd7tT7y4MD5/R3wXq90OZiVKId
FCB1uP5TIFcvtsYkIglflCowXkk4ZJvE99DHs7pqCb/wD+1We0C5KKDlqlcjf0tW
XjeBtqzSu3MynRGbTm2H59Xx8nP2jsugLuM3bFkp2ZAsgX5cEK47iEY83fj6vIWR
OcwdjTseHwP9ypQTLpIQ5ETn0rnjRgLwDalOxqE35T4W34eTkQ3XuMKwgQEEs2fk
xvrm0s2NNJB/3vSdkqY4sm1zX+XglgP+rvcywAWJItqL87ZLK3m3ZG/pY9Wdaq+c
IeVdPTfOZQKdVVmEyqUZ+rglfw7fqhbsQp/y70LWHRr6fjahq4fXK78HZEC1Bf+P
slftIZk5hCtHO8k22mMOHHcmUGmEobowtPm3sq55XEvOqFapPGi7SaZpZFJ0Bx/0
Rtqoy/VP7F4rjQEbdJ5uXWM6rMEkuyJtPsXYiqM5CwBw0TOVLCT5O4Ie7zhZzfq/
LEqJWW6eYHE+v8MLP6+JMcRFa59GIYuak86E+mWfIaRgmhxzPeZ0IuvvkRb3/7Fn
sDiGk6OZHSTUPQfT0cQIh3Vqth1fBuS2a2AW+LrZ6oMTm7ID/o7CgCvi99PaSZQf
Bc5Mzlj+rhK1DQoJrj7q0DliHK0ZudwcMydiX34tU/YrQ7tMvTLWRPoOPgDbYPt+
kJqRkYlX/m+AcbHCvvN+7TwUN/oYgDG2JMGV0nFEaSdBrQfyN/d96Jo0KzH7PZaK
Xlm5zRdu5vhUP4KmZukp8veYmVXzSKjy9gnpp0ZsWttAJAr00kKB2eW8t9gmu7Ux
s/3YiHA11EGKwp0vsioVdMMDPqUwLmsz68YHTckVIx0aQcySacMvW2X/vt5Afgdt
v+SmWHRqmPRNy5kmNwujhZ/iFJslkPiZno1NPkMJGA+Hx8q5gAeLDsojGERF+0G5
Y/tqhmDZ5tOFxssekzEx+rv/2CqlG2m8XsbgysivVFHxb/a48J3yO12jbMsVfp82
4ZDxg2b5/CXhoGXZJqiO7jXosbN7FQ3E8DPFkjzCRVJ64npDbxo5S3PBm5Q4e8tn
EJoL4JKsSX4CSeNZA0qY7hCt5fDU+qXPe5hWzGd2clRGO3BCs3yneX+G9nUJa1CL
7H75RkKfDUvEbAWO+cGv0uDp3setnNeeyxvssa3+GfgAWpRvirkwZXWPjHd7f+Nz
RW4vIOMdeO4ku4yEPukgXICeP4vyJwgtcfRWuD6korJPM1vvSIH6AlEkEgufxY2m
PzYG5Su3lhgVEvCiHbWcKD1AFtQg0dRIXNA+m1qaDy5wkvtnZ1snbO2hqiulUmb1
TeYXkrSJKD1H1skMm7G7DMZz+jcxyzZkEUGaM5Kw+Nnw52Z2cYlDdPO6dlz+trXz
or7xAtpoZfKbmGcu71aCB3fQjJSYT0XHu3sdwOfRU8+w7S5ONy8CkES0/Zb/8NhO
9OUDpuChLskK8MwCKDMB9mSVImkOdDXzIyIGcEFnuR+DHMjLBBLCYU2EJm1bxuAG
ZHRI1GLX6r/T0eH5+1YTQV/1KxZq79VaSlD0df7fOAhRHK4Ic5CiACMTLj71ll45
la7D7OXUJuJg5k4mkCGF7vr5Dfl6M77fHAMySiziMIQP9y16GDB2B4cMv0l9tqBj
UNSZQSveL4Efbh0vSMjzsAb2RbmQXEfymo/nk/iBeiuREqnGw/T/d/u62t+KAfPE
cH28xPyslZxUngjxM0+K9ORcQv5/lhPKReJV+IOJXpdIVpPX0YkgW2LI/DvUlQru
VkykNLog4p/XdDusBaJ56qoxAQ3BeMyE3j3GbsUWiY9ErT3bSU/Gagip7u2QnPfM
DdBYZdihcg/bzBfS3eFFs7CVUvaQ74sdVIttr8TIRx/BHEhPDJxOSwS0XCPLP8KE
VMVavoIWQiMfg/i9sNRA1edJdbQgnNvAqxLfGKjFXsH0WRx9c2SoFbYGwcswVnv+
Rh+4/o1LTNwz3RNy6c1qZX573k/et3Nu04UDzUFCAJwY41ENWY6zVTS3pOghCmLX
1n4TPR6qDc/xJSUqxXO5cbHBr4pPn+4JHiFXdD7gthu00i8bNj2FVnQMVPUmw6JP
NFVhwu0iqM04WqS/t9vOrwO7EIcFytf96qJlgnG78JY0Pr5KhwSvRfY47jeqFzea
Db53dHXbmIOPxNaLXKjN1t41mU2fDmF3lXGqASOPP/nis2dIej3LgmFZc4sEzPdd
MEkQDns/pDECX8ltUiq1MzhZBpd0q1qkkTZGTR+oO6mnUbvJ0ynMYAGl5877KoKo
CwPx/bTD166O5TbscsFsFGSK+9FjUOID4I5L+Fc3L/IxW6KeLOBBsXPXXwO/aF60
we0gITYRqfvOMLalDvxQE+YJ6Anne7OWeb9HIHLOQNHbY6KATR6vQ/mFQ8n0gOwC
H+giMrUXY08d8sxjgOD584ThOPWLMCEGBbQjjTNd6ztRomA3bY1eDVxTxoS7kXTt
RJAp1dqC4/dLpaFiAlh9kO7tDr8UsHXMDciLB48XyVFU7SrmiKIw2qEX/jSlN8mj
/9gEMuYDRuBvXTJoIOtCu/z26L1Ms5rJuC2ssfaUka7xkk3qRmxBuaRnY/c85n01
FAtBiPoqqB7zmgK2Cfm0CnAbA8EwT1AhHuT3So0kpycRCEKv7swxjQcuupDfN3VG
BFtVmztq+AHijrp4UjnSk1X5IfboExdTfC/WXhtwRyEwV1LGeE6DE7Jl1eK/Fcbg
H0rKp4bhuCAgoAxm6NqnIz0l7RYenyNKbGj6r69wDIKw9cOe8StL+mua8kmHyHRX
ppofl+9PhwloK26oHEWPQECkeynrK8il+ShPrIb94cKrz0NMLbrG5C85SBchqzrV
NjSO2aI02Hr65+dTup5NAHrikjjHa6/Ww1HVxc3OhUs9t6fVTbCbW9rAc/vt4Qj9
RifQ9N9dfE30wtbHp5/5gw7OHRu4BGjwQVssDK9xRgrvqfnzu55xNb/YcXsYDWpr
c2rGFLLbevO1usmTRmm189n9Z3gEkREacOmhSbLOdV6GwZ2FE0NYP4ZNdoue5Bli
NaOtylWg/uU/tAovTtjI5dhO7It9NSY+KhDDMuLxCF2LLT4i88H19lg8h9kpp/1w
cy8hnjEjCwwFfQkjI1A8WTnVDFx/NYEFv7wPWwrTePcm95l9NdvgJf3IHOkMqqPz
UozvIN7PzjBTEd+5XEn8XseeHADqx5UFoOOaCp8/Lkt/V/90g7asI4bn2ROZBYMD
zLBLevZ96It+gx20+RbvZXH4LXA2Ye1jGnpgaotXshqUxok8/bA0P1/Dv5hi+lVA
l4hQbwYhlKTZH+eGZ3OExehq5/IeruSwllXZrGhOWFJR6WAONakCKrRQEYowEyFG
hckFWXZKhlEiEvvpGQEIsIsBygTNMEcmYMafCgW0N85OxNCy5ChOVfxbHBaUDMhn
f8nnkFWg7HplcuTxjrXT/WSeqlBMGE9hDUI0C7i/j0upBxdhd1kkaI6byjy7hWp6
LnIp/UAJpbtecVcpO3w4sEicmJpzQXvQTsrQp6zwmtbT2juGRIbFgNARuJNTb+zj
2xuzwtGBFSrExW3bFZ7ah4muptaNmYxsZMT+FZVusPU485+dtgQq8zoeBa51sNOw
nypYdjAOXRe3iEDd9rU5TSAAX5JVfUOkR/ALPoPN1dP0qYAfJwDGImBoNrTCjYJI
NgM80sCPu/zpEzMIMy8YuWzH9W+Xt66l8vbiUJSLvDA8bjyU+LzVvTPS2vw5Bl2p
YlW2rCtEIOQxxpHP0w1Ary9y3BgVr162M4Z/29jUM7bRP9V2lHxYU4RamXl6xXGA
q7krJFEIy//sONp5+PdQM+oeSHTsWiZCU+JP1naQBde6XikMjSw8WPTtrHM/7dVK
aaJPUhPin7K2tfwHacgscJRSxLGvd2UgPwGq5koIrfdU1Wgzn48DR+z86iB/RG5w
o9z6eGTt+Q3ieWBoT0lhHQAIY2O1wt/xUT27iTgsqil4Kz31VQjH9uazR3JxpSxY
RS3y/n3wMghCAiujFHJKQ+8YFSTLYZEhzCmBqatEaE1TsARLhTtCrsbhaU4a6WjS
Cln6q+9Ol1TsfDdnohob3E3qOJPeo8zefs+bHWtf1lBQm9Kw8STUBQEOiyqkdJFT
6WhR6szQvy839kL7jt1dg3ECI7Szc1O8YZH2ybNtdfRZNnKxC4DTcV8sAJi6nL7c
Dr+2k0pl3koPogz3DYP81kOxSwNTHHc116q1z7YeSi9pWUcr3CTeMtz1Dt5qSXpD
Eg9X6CE+BK09p6AW7c4PR7IcM0vPEOonCmJ8EWsSHzOU20yzfr7YKZiHLmBd9d3i
jeuHPxi6uiZRpLGRcqsaBDNBeFA+HeivjmbRaX+N7gqLp9GcZomodZnYWxo5GHpf
o0KS7L/ScPjuz6pxKcuDkISn5WTZ74BwQOaedrUu3riNdzsD8gOls3MZLjgK6K4r
nALRL0/WOVG0ozky+cub8Fpj1zxOYrUNU894siIk+VnSqYgHN5hpJzdgjDlYWPvt
nLuZudbgj8iL9T5z3fOrlw4HSv60FuhrWiQQVhwgebCciPYDtricnp59dNfKn1fb
7U8hCsPI95A53kRLJ/ANL/K8JjoCAnU4xARcJdg6d7DP4PJynUtTsr9fidBc6Ura
dhv59bm1loTSZhg2xq0l0ddyeD/u9l985HnDYgaYUAX6usRGQFvdVR6knFkQVkSc
1u6nZ+7/CADC5dAtHTb9tmyiZBeM/4UxKvasS07CrLVZfFv1e+7Goyyb8/D8nkYR
c/mIUoeH+8hPxBTnph+E5Plclh4WhhrLHjRfC/CVT7rCchw7npXSoPD2qPbSN3DF
0UKmy2H8PNxpLqo9ToKyQRY2EwXYtZrrwq7WYGkWG3twpWcs+TYgaD2C1MmuKp4n
vhfMk3WFXFiiHlMPpojHhXljM8MlS07yaqRqTHX978vG/GgQatI6PaSo55GMGNNs
hxnX6ZRL6+ZzrgqDzzeUo4GzbhBIB4SBijyGOuBezOE92Tj6sslZ5PzCx9LZjNtH
dkVe5vXaihFJ1F3FIT+FcF6CkzIyFtXAVoi+gEvC0AghpW5KWlYuF+mSxeM65eIa
h+aieq6RYuSuPjnSRnP6cItrRxrig5WEGAHbUjb41mW/khUKJBQxatq6Cj5UeZ9l
rhZ8+cyz1+Pn2OkBFl/dQys/cVsz12Y4V922hiFL8b/2xqzkYYmBKwIvuwWjUtgw
U9d4GvFr8ZZo567nCKinmxFm/K9bo7f8JYVEdB8F4h0Zksyg8MQWmu+nfh2n7OSN
CPOcRZdiEOyBBVm5oZlU8ulgQXsaE34AmkMmMYZIMBI+fpNvO8iYevhqJDkFOAOa
/uLNEjQs3eW8LRGmvijRBmnPAYxJKrHa3E2nO7emEiIRbewD/voc4MZlWuxi42WD
K2uOesYsX2kZHU3FTsCoTIhjlHnrJj89kgbTdeqdMMtsT6R7YXvTlhxFZiWQbGmv
ZT49Nx3AQ3jhJg5xHJoSsipM6vyhqw8mobiaZMhqMevoh4anXCzwX5zk+FlEnWGh
rCdR94fBc8wqUHIyESQpF0v1lp+hRrA1obHS8yhInAsTbZd3QEDgxvPGPmO3KWrO
nxdaEZIvkl3CM9fKPRN8qQFhwa5D3i5xrmvQ8daSgWz0muek/q1BMWvvCmDtFnUj
w1elmf47hPnHN2Ood4YrfLYQu0Up95CEMcrfiGsoBqHLtFxieH8wBzarBwNpv7sc
U5WLQpDxN8v1vPSHGwGWWMG1+3/H6My731hmXrG/2bpFdaZk7T1DprvL/qWB8SUS
8JZHEDioJpuSLIEoeLT8k5W6qKiu+f3amE4jfl0Ovxgrkl4H1LcX60Ol7M7gCyk/
LkipQ2xOOAXHX81frWmFP4tc8gdjFg3q883aSDDkcp7SKuwCPwdxmq1E8EBtmMDM
Kis63z84DOoclg7Hm+p32XMfZiaO+Vuxn4zb8yPQSMCAyC6tx4/Mecky3jLVD44K
9jtNT+u7z8TLKsIGV6FaSoD0MNRAAE8L/Qa4yddQx9dcseIKdSP2cg2wafZDy8FQ
PIrYkOoBHSSI4s3ulUBEIJvoCFnEB83NujQJKAVxJRflJYZHIK6w8xrA1APo32Oe
RbgoqDtcF1yp8O6GwsrhOVKYkXjmLGZMhrNPiLzRaoZ0sNiQMs0lHtu3qX6zvxBH
Fys7Razx3eNnbPhww+rRpxaCmENABG7ODpL6GED/nWTPqcrCsD/IoZWeOpO3U2uz
jjhRz2xtwW4TUKWDFmvC9a3sdRcZ+XedCU74m6cI6X/V5+3sHAJhgffF2JlsCNOd
f4X3MTkZdSAjstLUdIeAEqwbuTaC4LXXN77YskKxZAJPhAA1gnjxer+6Wm0v7otN
Vl1fjYffXqG4h2IOuqkqfMs6sWzKy5V8YfcGD02+k1nUu21hN+6G2SPWeAhwahPQ
4ML6TkkZ6cR/5O9vdL/vaYdBKENSv15KzO/bu7b60YVmfEZ2Cv3TvBeMMxhWFU7R
DoKS9eAZXe5UfUt5qvGMYfWCRcNJ4fkzp/UeI2O1qCth8bnm7J4sLx57oo37mKz/
28YEMMZ89aG//+WPDxfL5eLaUf5LUdhCE/W+wwV5k5fmoJ0B7XHuFCQBOWnS5wEE
Ocg46iYlq2P+QYJ1w4kQNSA+bX2ncu/R75FY5KbU0JlADwfIwuKKPr2iyuAfezoP
x5TGzN/4ZvyyCcsnVh4mWZG6jUKGkG5LFJND9R+md0oiAwE9AZIdZGOxPKAhhkEs
QLVlt/041H/PknS+gB8RxQPwvtflgOckvv85o9uprjxc58uyYdwT0OYjvfMJYn4R
AOn7WxRCeD8KYtrE3PimCbCIlzSnfSCnABuRdsThkWkCb+RVQXq3uxq3UETxNf0A
D5bWP/Il+en1wvyED8ie8QRGLnolNBkFk4F6hSoj8NXmnqLbre131/+j5gUSk2Mf
lZr3pcv6E5t1v5XVKAmNionlO4NWxBc5myoYyae6mPa11vC6RjaMwvaq67W23FrJ
6F5YLVTHprnY/zy2jf5Mq0qfvipYrCtNPfmvVJi+HjDd/XIwMynSxOLxR2CdYb74
SruA18oK7YqLFiys/eNHzfiwgLlKjtpFM6zHePQLeJS0i5PJx5wpn4bob8gk9xLE
HcjqI9Ixy7Z9nQGw61mLeO25anysashW2zaLmh9pfcbtEdETKrkE5jlv3/e8vwd6
TI6nfXNwQ40myxUtAqugtulfl90sHI4x81VeyE8bqhEfTdfKNrIxm6bVb3oNxPN8
SK/bVMqrkL3FKoo3+268WxFMJVQ5kv2g9M8MYYmsYdeOBAYCpd/F+piFLU9+rF3H
Vggly4xVk2uU7RelGJANNQG/6io1ksexVKe0y3BtSfcliVGkz4C1ZdwRix8me4It
yaI1VmWeurU2WE6mhrSkTgLlaXT7SjBkR5vXqNxU1CE8CyNhaIbNJMy2Yw+XlTfd
ugMpT7SxphgC3TQtTEI9KxP+NNSXXzDbTQwJZcPCEmPJWo13rI8BhQMyFJsIUHIq
cNAwMB8652iTb1cc9GplAI3ltvRDzI0Gk8WVBJpe//RMM8aMrRliYbWdxdWLvoDf
3lzMo6+yZrsN6kFClaJOhdl3UFLrAzjbD9BurEXQfyEsgZTxYEdMw5PVgCFmmLje
gy8KCskOEHK8mjsNjltDeSc3QeSM2arkUrDNeXU8MqqenkLcZN1BnZ0c1eDMW37y
7xHApHIrFUy7gJ3og8sfaOjQtHzXKNXaj2jXT8JIf1CBzhKVyV3JQH03Zc+QRNza
NoczX8v30nNX0cfjU2ILSm5fDprKNlosuqcLfEl/rQq9JpZgj3CssQLFAObYnva1
zRd3PWX3l9ZvKbtxGop1Gi1myzBxwx13zSYKmAgxJP8o9XhGcvDZos3PHdJt+FQ3
Jvg4QqQ2CbE52ok6mkVGOLB3rlSWHn0P0UQfeJDj6Qa7AElH9+JO9JTBd05tTEdW
dAEIm1xngxUtGBv6H22UxUhcEGsZY/1Zj4dXZ8nzgGQbTVEWKZBGPRTx3VKl9XEs
Lzo5EhNA4jaWKfgQiDOrqrG0n1BJbL84fdA3adlZ0p5jLWbilEPSQ7wH6Bytlo+4
HbamM4Oyb5alcep6IVLmo5t7ByHnY5J9ISkLDciJiB5HuttMcFHaYBgUvh+DrT2Y
KEoLlXgEWTNWD9aukgXZc/bIfF0k6MwmRjavyD6dgDL8R0FJ+wUuCX4pTj39vtR/
YU810v436rzUQl/kDAie7DZ3V1Clr7Oe2CHjsI49QsXh4Pum1xbXvrb2psp1ur5L
KR09CuMIwhNve9g0sd0V5HfSjs2DjdqRh/fPTNOt/287MpKdKemsMH78668eJiPn
kPyzAgiryaivaNhiqBzhpOZ3EWKOPTk031mViVC0649UMzuwoOv2dqseUwEJMt3u
lD1/Hd/tg24e6Oug9spfL/xnJ3ZzCH3QarVd8ZMC+tZtWdBZrTro9boa0ZV8W1XT
2uMvNrSajfqkacE9U1mJ7O6EcHTW6959JPNYfMA9AA1v+7EamMy/02qB04ad0C9z
+HxTj4qBEm4+Id9pDwErBUQCmyNa0JZbnp5W7Lyib5zBn0AMbASwucLSBGG2g5KU
36KAz8XIhrcXivin/Tu/hZgIEpPZcJ4aarNWHfoledfpNK3+TCgeuWv7GTn/YgPH
pQS32ZwKsjvRN9CB76pCus3VyiPil3UOkGwYyUVF398MeiglRpog+b7E7JLvvcMD
dR0nbPjstJyUShuWPZBPcgYXdz7pwshI03OWSKwsq1SDU22AfRyE9t1cXj6hYLzv
cbPHAU3hDNyCeRpzKjbQ1V3TuT/JidpD+wXVU9RperwQ6QVuR49c+p++3RPx7MDe
Td1Gwh+WamVb0SF6i14kJ3nAXfb0bFtZ+wm/+nA6zzECgIan0rfnt4/jZZ7AW80c
mFMsiX1fMK+pfAJDp5zOy/KHfg8QrN5A1A7yT2R+6+v2dyTM3X9hG1yd5/UdO8Rh
u3eJb/MTjLTd9ChNDIRiToCE5GTHPSYc5GkhwJyM+k0JYnlrT2CASFbaAGokp9mH
xDKvlzYIk8yY8ciMLL9qy6E9ctwjnhnoFLv2VfCylIlADeS8SbJ48EUgOuvd7CDj
GJY4CHszHW/DsDkoKyaJRqglX9jr+P3c/flDvGdEuznwURe1xkAwm4jabPRYlPLd
Yt73TuAsK6pz8+Q0GNDLI7inWQodjh4YAF9CW0k/4+JFoWqYnge0ixpJ0whf5JXA
wqa31uWHiZShFDzcnlbt0LhzQmGn7i2lTbTJA6D1QGzuWSvwcn7dpe6P1Iudll9E
rz1ScEMQM76HTq1ZodNMoFb50IE3tssZE1gnXClugQIT9QMpVoUUA4BapJ9ASSyP
3QD2NCyHZfOwNqyd/QfhH3Rjm/ZgcIGllzsiLLC4O6SG5JNl7opDi062QdZJPLLd
PMcIMJ9ZChjbNet1erKUyzqirZHh+7J0ZZ7nkhLFiXwofeHS+xyqrP/WH/uSkNxI
b1lngroSlSrEFQhkeZC5+YmH3GCj8VXfGXp4IkSY2o87toOuVZSOJn78p7mbk9qw
1t9PA/jFe7F/3XWkd+VG9QomKrwDLlhlM09+0hlj5DQQUlttnOBlOOxkGbjhwQlY
GgHBy9hXVCoCIC7+uXY4bWQwTTjVgQc4xeyB69L0rqk2USKAqk1v25a+HnGAVTVj
yabumL8P1oYXuBd3txwpdhUs0LDEDdnq/SNCpXj5yOoOKet7JcQ3zSTsW/4YEflR
Ams8Uv0ctbWDuD8K0n70/JSkIp5umwUZJlWJ1wWwsHStgu1Q5kc8kRszM2hl0B39
v0l+IQwYk2k9Xd/e9LL+WRjazUmgczHna4cXzEsuWAa4LGfWOXlOin8lVT7tG8s1
RaoJHqq4lyn/PNa3+y/JWU1PKvMkSX5GN5sHVVNTFk4OiHEwhd3LaPLSbCLvo9Cl
n4InPNw3teehSfZ4fwPFtKoYExZ6Kp4/UiPDSM3W2VW/Lcj/3lHNc3eC6XxMdJiw
dgEr4Pl91BHyGk8O8owxgGqJ69Fx6q+JrDZFhCte7Dsz6zccj/YyrByIVbr4ra30
woVZ9MyX4OrARiTGmadDCubyqnG78AfjPIhGw7AupCmi2+wHPnQcDr1Iq9hLYnD2
5gxuED0J1uflg24IWMbWUHuqr8zQF9UqShj8PdDZKIKsTu4N5k8qq/cmSuJclbwl
viliMPLfNDqwdtaK41OKkVRoV9bsYmrqh41g6jsY+O+W0f62wY4b9T2aqwzZ6fwQ
Lf8Kg4FJCr9i7tPg+sl5ABhehilZ/d01nYLA51bjSfnypQxDYdNgyRhmtEYqXpSb
xCl/IPtCs0nSkkNv5MDIg7+sfcDTH8oUAxs0hT7mZdYh2bimkzwBo7W3PxwbBTmE
Ds3h76f11K58y9jqAVJb2PzIB2BHBCAsSuJ2sPHCEpTlcCKyjhFz+Mk8ucVN3Rjf
BHFIL3j2l6T3KGibheLFgeRO4fF2ccycsVhCyqA1hs/KZy5NctxnJySbZedhN03X
hC5cjFLP/cDOSsBRxD9lc4mk5OVnRkWudrjKVSc3NVEhhqQi1ue/4DRTOc86Aw9N
4pgPBwt0gauEhIO8YJNeKm4SjjN+/Nx6D/lm0gC3OGeV4q//byD3MFNhLVmqmzDF
GX4bcPmHWBgTDguncC9PONMYxRrbcnaBsahgV77n8dSA1Pfhgx5OB58cHYeNKu3N
pvgrV+HU6BGn4J7YVzv77MbbD6BPVA4z66S3vFL+lRQgJBlAcVKtktJrKtvUVUcP
0Rleb0HLN3aYMp4nTPGWxA/QBa9n50oqSEAcf/APgLSZec6NcCzbpcY9Et4Q9tFv
wvR8h4AoRGThIrRUPN1n5IiiE5qeaLq8CaWn1avxb7hiko3wly3YROgHO6KrMvMf
uF5/sWIhIjVYbpbl+huYFNAXPlFVAx6afSy7lQM0lsDBqJZ3wf6YwZMMNdEzY9Lu
0N1AIFIT/8saiIH18VRBlFSfg05Kaah+oxDWyhwy3thprB5cPXufEZkJWqu1UsZt
Lf6DVa83McAbV09ATVW8Bc8K/ISq+tmDjhjk/pLhPIWcbU8KzUPM+NtJ3V1vaIVT
FIOd8cTMCSt+3UzENPiygLkEpdranjDUgLxUX4TP5vHzFzX8tsiALkEgyqmW5ILL
iuLRF+UU/i6NsIXAVrqxnwzVD8j0xnKDeUzkzcEex/OObXb0UwREfPb2OsVEi5QT
7jN4qkL9LRZzM5tuFBhiwVdGusn+J1qoRMuPXxdDdZe40UFwAcXRsVH6qgKFZcL9
GjAQbI2SXPgOiYsu5ZiZ0hTQ6N2tJggdSJnvQE0iN//8J6fZ/lk5poR70qr1KF6H
zoko2PQ4KWRsYnLzCDMsn3h8W8EtoFetZaFma6COt9O4Eeop64TnVt/3JZOTj/sA
VgJHYgyR2WcPKilTGEuKLp4DYisgFjo36wcCNd1QE0MFE/iXgRqCW/JbnDj2EGxT
vwOXV3RgcQC1cSoIAnBM4oDnuNts3qbj5oZYPZ+P8y7JbG3SXsE/GfmHyx/BA7xs
efAfEtvSid1kfrxkNnQqrYXMGtYMDr6hZbVdzfFyv3qLK18NTKYWdB9rkJu3jpuF
31W+TzDCdW6l9Mkth1HIx/F1IHdawMfvQm+y6tp/yO+4zNrYPCZBvDBeiHsIFyLg
Hd6EZFSqrD3GS3WweXTNHy3nNysag5rAtGr2aH8kC5hGv6qUPGjsEkkZLcuQOaYi
JSNujqooVtcoLm8iZj06nAJPWBQ0tEwx7GlfGKS9A8xN47nkFzMI1BsUjWbe0lEd
nnzmZNg9iepPKIBez/bha0Fxd0il6nbwGxnxFjavpQBmcVgdfiiwahG9c7sXcBr3
KWow4N/mLmA7rkSGwGZxcORbuLcCS1K6Hd5uowcsHdLdppZCc0UY9InISlXb/Yg3
KYmlYOCK5AtUh8nCg+3ieEBolJYl5lvQXoFkXf8KpAaz9SBMA++weFfn3INhCSpa
eigOXDB3rD/EqA95KP9kInZF6QTZo9uwvcttyJ3BatR5KXaV1ZeAQFMqHQ6Oa8VF
pCESZI8tmc3S02jHDIhnTbK/0r67+/ItGkUCtf8Hq8y53NfMP0ioqnFusM6wdVDx
AywPzGXLAdXR6MWijget/M7qQQ0avmiTSQMFL6s2Tsh9yThiFa0MxR7NQB58q0ys
TPV3SVqJhK6NcZXNG95e4C4YyTc8kICPekeSiE7w0PA7r+sdlBEgL4zQiDlby31W
Uys7WACs5DfSmO2WLCbGTZr/g55pQY8e1KzfSFQx6YD34bAchhk06ZITpeKn/2qc
z8gZJIYWrbhr/XN8MTC1+6UdA86u69U3tU9q2mdvPYEAkDjjKyBzROHHYr9ecmVX
ZbHPcis26z8pDsMjo0yN0tWv/g7PS2C6uxW0lhwUCb+4axrWVKZtVu7bHPcfNpH1
XQnUR2CSWGL6+/PaYTQmX8sMwVKHjIUFaAXzdiiITCzD84t8mwGLIIjB0+K0ofPI
JAhBEHG9eEjjMY5MbsgR0wh+/HkRHeT8B1n6JOD93lVCSXp8WZvwogrKPeT8GmNj
0u+NdM/suT/f8/KfITUouxXGsKkWM3F4GmW5ffABugJb3X28qjyLX5Li8QNAdXMh
IL250ONyIBNIVa1B4qiKW0iCa9E3/Lqf200iRIvSQPZktW8xz4qc6IfZqLX3Za43
KPjDtOjmRikrGybUpu5nKbOuyrGrlR4q3bsPvb1CcV8=
`pragma protect end_protected
