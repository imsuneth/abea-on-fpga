// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:04 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aqjXjbfmj4juOrMXibopQR034HYe5lwv0+7WpNdxaL44iv20lDH/RPFvBoMhqrDC
e0UwTs3Ft5pqvgZPPeIMtXIz8jrwgX95ynC2NyrCKkTygi1X7I00ydj2T5TtPrJo
HujNYhyCHk65AD2Rqh4kT4U784xnHJyCq3q22J0N7mM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31664)
69hyLDzskrsXAdUCuAbPJEZ9xEGCqJ8K7tEAY8gp0ZF+MfKxrvJMs3Pp0zI2Nny0
2KkO4pt/kJp3yByzXtkUVv3OZDQ6tpjkKsflnA/F8Hv+qfDy/ZE5gf2gqvREJkbA
6OW6dGOumXogMap0rnot9xKZY4RydianhJjZrnIwqQ7lL2a4Nvu5LgtKN01wtXku
gErp4orLoGwVIjZ/Yz6XpRATcNqJTA/QW0ZSDb0K9581alDVmgLsZO25YDRGNmpt
qKUJhHi1u0wdN7EJdmdjUXWd+srMSyvIi3v22NdEV0wh9Fv17CMlVF0rdNa1ZLkr
UIxXdF9ybvHxeUtg2tmt1zWGveJWE/cfTFzfWyYzqk0gnOrsVi9wkyPFXynSZF9l
KJGqy4W2LbzywjjBKsOYA0C6kl23X2XdagIbo4Mb/GcNbZnYIyl8UogUdFT6kLu/
yYp/STpyBfI7c9Xo0AaJsbu2iHoHloHWOjJcv4EJGN+XSDVyehM52QLTQVyG2Vfb
2PBv6o792N467cAIAAz7Mv9aRxmWREZbaBIKrbLkLXOaY88A+S4LXRqmbzqYnn68
Ug1Bg4GtAcII5t4pagEZDwRRNt+1X1OXPrFcsGMqnJ9Kn4Q07q1Sh9Y+w5Re8rNV
ssM8917p7nHc1oNHozp4rUyThOLxjnOwLFbX4/ZE2Kiqw0BEbPqQv9iqwMVb8RRp
SVhBApTcE94sDair2xsfS2K3Sh7LjlnP1uoOcpseiAX+tgS89YU1RZNsjSOQf/p0
BseIcft2c6dmpgeHTTy9LhdazHcYchiAtur4OLP7aFTy/ZDlXFCczdOjzLLvrjUz
cD/qKYabnebQZNkYjOMYWSuPO4hbw6oRKiPCLozQQpqbMooLamgXPmyZstqJXLP+
QMdBbec8n1P0NydLDx6txhrIOYOqYTfQzLAutCYik+7IGMPlX86awa79qGlzS+zA
s1dEwfdVqaRTAj+DX0H/LIY2iwTJvE3fvs7iqzzH/WHk4LVB32QKUe1tFg8yZSup
0Gece/jtjaoSG/+oL8xVKaRs6Pd/gYRZurNNpmHDgGnU0UyfdXxYTzbrQnmUjoAM
vDH+PQEJFGfYWSjnCbEYgPd9MNOUIygNKY5+PYTtx2emuLKHW+JVoTqK8Dv9Is13
wdTgnRC39UVE35uZquA2gfDwNN57BKrhyzXYk5aIyT90QiOETRWZwuPUFadk2vFL
3MlSH/Ca7UmW8OwM33gLchCTBoB6I01B7bi/MI7VtM8w65/xC/AqaAcp9H8xzebr
TedhmJ2CGivbq0daTJJ1eCPb20cJliNrHOBhCg6rLiy9Ghw/zWArdHJJx8hEirEY
L0PJgww1U8Vl7AzrL6Q0rqYqX58q6oBMY4DWhhcvL9B9sVU76HVS+kBSmeP9RlU4
OYSn5pteV7yUi8ZMa75AulI0aMU68Jw0yby/Ixa1+Vv6tXMSiiSkcr5bHiQR94J6
aVsk0jqC844XvOKWV6PO9Wx6VIKTzKAnyaEZhX6893zYxQe1f7UnkQ4uCfobDM1n
A7ZqSVZKCQ0LmbOVP0uMNXKP+ZdV4TS2swj+x7oZXpGh/8p3znGM7db1VrRlmEZV
ayCKrr9h36+ZC1nUOmOwRYEfCBxxPWOiAmWyBX+HW6buZhDitJBulpNu4bqJFKiv
Us10EjGU9EFxF01AvGaktmV/AKa7rzHJbZSY4xK57+TRFz0JizUaNDD3H7dbgF5g
mPhHgStgK5G4zhu87emog+WZ1RXUGEu8xg3yK+b74i6+8wSauhtEJFHXIkquQwAa
tK+gHwZt3REgkv4luVI5hDsxe4JNa7CxGliFU8laPBQZiWo6FQ4iVuIXOmOVJg30
3DGbpwyrctfrBckR0XvTL3PqoEgyLrF0rsGQAWIeeUK6Ke0wE8+s44YxrYRSG3sG
rCFy28KP8eed9XTiI17lfRvFnsrhk6TNjpeP0KOAcgpz6nVQEziAqGolM4PibBPV
pQ/h8B2zZKIB9XV7m8ovWTbM5vpDIrwSumYi373LL3TiDWtqhXJklen7zrrFAMWS
Q3dUKgVRki/mtwtXSWIbgkTzxqmZGZzyMXIk15fnEdGEUggm3VB59dRnwPRmmvLE
kTCVVJFm4oL84cyXih/6H2fBYPSSW0zKIEIZSMLY0frLwNNAtc89sL0EA84dMyfJ
Gtr16POS0nNpecnpuMiUS6Ryql1xku2SeQ/2mgGKMMOoUe0IaoCrQ8eYglTCrL61
4BvkV6bwIg7MQelVlYOiRoLu5Q3ff6KqxRH96ZeknuVPsNAWpX3d/43onLUvfbdV
ETcWLbPHL/bx9DW9Bh6Ex8tXBSl+7j59b9XnoGVVsEeYs58wP2n+CkCeP9+cHF0g
qwOu5rGqXkmYWGQfpRCnNhpmyD4lFPCDbGXD0/CGFUhKI6BYezfHno/zc3oyMiQ9
1yiPhhAy4UhZSKKIsTxl39Mhz2x7RiPsOS6AtOdcqSaiWEqJE0cVm8pZa8KPzVHN
DkH4elA8Wr9TJsBr3ynjG1XPV9VSQYq/4a32XIEgQhSAQq0tbNsSFqD+On83NcXN
P0Jl0N3E9XSJnjvKWBoBEsZ70W6egp10RDRxhmr8x1yUYGGnmuqwvZ0/WjB2skWb
Ld7kjj1AWxfRjR/RBjEQMUFJtjNjDOXKTMeLsvrSJYPnNU/woUteHVwXVphgOd5I
G+iFlOMIgg4l8VwKyfwHG7fcSYG8jmszDkKEy4+OkqtTqtIdJ4WMZgxH6FQSax3p
F95tIeqBidEd7MlJThSyqE8wQxywGp8sOHL4TiL1t7zPkP0BFQWYFfWQSsQTzS4X
E8aPL4+VDRDhLSACwdLM+Qf9AKignOoquMdsqxRvTYOKSbQpA0XnJx4mmArAF9Fd
oBqlNa4Msxqcc4EKtLyN608uctWokql+G2UkyKM3htaE9WUeOgf6Q176FUCREbLC
5CVfP0sKQ3s1XmN0sSaS+CoTFmKgU8D8J81AXmtv2A6k0FEXuSNaIdqx9EKmEasZ
8GAxapFtu11hDBoQQW9FONPt7X2CFZLXpFZ5WX1Vty4AKyQR0cxkiDxUHMNUeRuU
YPdIKzyvRaln/RCo5oD86kgw7Zv4c/DbVN07ppCqQu7/KYJQpaaRbPu/85gBN7na
+PEMI1R0z8AV492lBd32TlQ383MMjnBbDsWJuNNixXfAxyEfoDiDjFBe/48JIt0C
MoFZXKZ6lAggJ59/8y/GzABR6KlkC0LWnonc0S+DJGocmuICugiZVTApjPbA0lVu
1fphNVxfjPZ+g3qs+DzNLJR+thPD8HrL2Rvn1n3/6b0hsFQItcKdGRI6liYkssBQ
yL9p/KTGnWFIJlrvgZmE9ov7EPYnrvycS5Tq3H2P6rtCWENFHOCUg3SovV083EM/
e9lJ5ORQb+otx/Eoa83R5GNY2HSOI5Ydb6xgc30HeQhoKgv+TeUGtEmQJ/JoRMQR
m2EPpQwungzOjPTfRkX+NO1TM4PFIQHipjxtcny+fa0wqlIHCVRCaI1URIpgKkAj
jB5jiP32h9QMNHgGu8gspHuVFUSGPGFDqs0VOCiUjnUcJpMw6/sDyQdhfDDcL+Cb
8t+BeBviuU1FCnREMDMfadktJzEYHocg+/4FwfwURNAA8TcLsuUMIGr+NHnpbfcC
+wmBe2VvSM1O2pKSxYLixTomBs3xBP2y5tN31HzxWwgFzgND6oMcxpFrV7gnNIt8
PRTKGWpnMUqQr+dakt6U0TdGgJyT4EfbEVEqPsuaO0B/ze78xT4WT3SuGdgKR7nW
wMSuLBsSVfWxGnSJ8iOFcQBA5bC/GCjS6iUiZnLffgoLv3j0Ra1anHopABcpGEkP
H7aIRtnMVbecz4/8tigKyLBwhyt5iVh5r+lr2FCtyVuudClp6gtPAaMb3KEiEIBW
nCVVdQyP0rRZ8ThXBWrUPMIb4nwM1raaroNQZwuGixSzTP11dJryzTCt97YJ1v2c
CrnyuwYKyL0tLmg6Bg7cJW84bC76MFrB/6hRnBFHebgMP0R/vPt7V2+suGE2YXz2
2XDC1seTAZWVc7QhajFAnJ5Y4n1M9dtwZK2B/YDtMgDhDgMkhwSnOBwzJqsU6fzO
p3/dIqI61bP9tqqrRL+81uG/5bX36Kl+uwx28eX1vI+Ab39rh36Fl6fgbha1iwGb
wNouuwmB17KVToNYnqk+GrkP0I3KHxTmSrfWxSAta+h83ovA5hb4d8q+GaeYcd24
+SM+v+x6gSqwsD86RmjeDK/hT46LnnOv1ji12+wpnYtH1JBhYUMShkVgpBOk2CJr
HQsT2FdXMCb8/tbHB6Hu9kCVnZFMKNBsioEbj+eM7B7UacS72Z0nWPwq9HEQisFN
NESwWSXYrbzXkgdKHTRWBDJw4gMyaHdAjbKxKm7xNWMRWUXHUmoV20G21r1b209j
hyAjlslTBZ9Fhfwb1hmhwTFYuIH6stFMizQKkQt6QVfasrfIJ0uFEXSvsjpLQsB2
/jxbAZuY2Skrf3CbmdY75woH437K4q03q7L3/rcj05AlRmeb8m81j9/BzmZ/2S37
TSrW/YUBqQkj1EJu7uwLZKir2aHtioklQbn0121VSqHb7k7dqlyf4jyK+Cm+cR45
iF64zaiN0GRsEU7lJdsWW4JwV3BaK6NHaoQMvBTVQoTcYHawlVl4WfdpYRbpp/Kq
fSYmZ354BJ4EuW8Tzvadel8Hqn4TcoCmaRJ5vufJyZW7Twabo8cXBQE35M3DAvmc
50Dp6i/2Q8IgTC/sVncnNx+QFdBEQOU+6E5cZ0ixWFjortCXmcZEaDY4jIL7eN+1
2jgsbztgInfWfuzyuRX4BoV9pxSQ6bh4DM7fKwHGzMdPiG67V/CXt4LhUiAzHsqj
0c19kEffn0ZsWQCKnSOxsSFvXrg6bYeJQZwP1okg5DMQA9cOwMpvsPIu0c1hKXVb
29pspAJulQ6zS0KK8bfa/hNaEcTQsB84KF1wKhl7BhPEm7QeqOucEifjK6tdg9Tn
MU3tQ/REAnUBuDYFC2l3V9ofmTp+dZtM8GG0U66fWTDJglDDk/Mw7H6glvdVKSny
gkYXO3fT2wdEOLoJD9RGRLQAGOrArTLXbyagvrytZkkeR2BeAmp1IKBBeqzKm/sT
Io1NoLy8Xn8ppHrgHe3ZA08wc3zIbi0h15CuTtDw1KZo5v1utVX5CM3QSNjcComr
CIAKVC0P0E8G6GPJm6UjBU3N5u+YTYQZz6Zu4/o2X59Z4RnoD7DX1a7gepV3b34v
nZ0AF0fhKyeelT+QVcJtSAxw1P2/1YUo146kxCPESdkIDJXBSkYv58sLk7koQLxE
qhpFnNO/XfJnyXhw4o4VEHpKYybJjlLMQ15F8g+Gut48bOmnFJCLmaeddIYhRSJX
uDl+0Mo0w6v1otAV/CwNpx8GQDi4vJdL9VcnDvLBUmgkO8d+S4/GZzB/T5oXN5cx
94zYnq56Xa8wi4bFniCP/U6cTcN4TeuYLIPoaDGZBuOXQE6vQt92NAplws+LqaUc
VurARHq/iinMQ9/niQCRRWC1zB8HemrJbU2EQ9fFNeYEpbw/9UUMmaDRCbc4h7p/
wnO5XYomDk5Wi8VIXwDO8YpYyzXbT7lgqzcrebHfpsG07CBDtdxVKpGSzHa+c5v+
1ozkeyqcveQzEVUy1KmdTcoiNKmyVkTogrGUs5Mr27ySwoCPQXndjEiv3YCzfSEI
j2YFOpi0XwKcLqDnrkx4uO46lnHuLLYRsZBIjlkKpDMLWWo5rUaaPDki5LNOOIv6
YWtuJNuU9nWdTMoSd3IGjoTR6bcsSW7E8u2OLq5Qk1wztyQjHAjV4rcuJBUl1qEK
qk/e0D8wLwtJ9KHDTWYr3l3OuLJI3rJ9/3UNkEHGPZ+0f1SrZlb0DsWcwae+fKSr
pBrBCvAGYjOkz02fnhP7HWDu7Gy913DIZCESDvvhxuhBmlB+ChXq19Q+CWFKcPbr
1L+VPIw+sdWhmCvtkoS8+1y5pgzwrO8nO+FcmlpCw1brmhOWEGxm5gRAMcG46gpr
SERnc7sHrjzCaV+yQ2LVLxPpLvz4Xh/qEZRQHothN91GHV8Obi3SxKdEjrdHS6/Y
I5XT8yEilWj4Z1rca0io2AkB0qVd37fZem2+1mWKDw3fekXwxJuJVuGP+fdiX1ye
9eYfC4t6tk1gSKjH8aEdnOeqqLfdwKjXs0fQlkhwBOlvcBsdoc34kHZBv93EwAVE
WPi019aeaCBCnw1ezH6HbG3kRYCquOkz0DzxJE34AzHoYe4z1k3RR1LrqfsQdjTh
e0BLo4QZY5eq3Mmu8Y0zAHdcAKVZu3prI3+IjUKK4JCUH7lbCHekqsDG16ZIsKuD
v2pbphLjA3TwckMSDAlusAQrnFde206DAkZdiBoBo5nmlsUbmT+boBQ+ftSrmDnO
vaIcSiyiwnq5uKzUzko0avQgwxKfSCWW94Bu1c+N25or5RwyaVOoH76DV92EnFwa
uWkYkJi6kA3gaUolhYXVRsHuLT5WdvNwFo4vUR7Plw/xLOQoRxI1AiRA2JX0ca4Z
lXKaWODv2m9c5Mn6JyRVAfaMdF8Jco+85WtbkWTmaXOYVzxMIujKlPdCgenX/JDN
z7+sJVrDbyHPDX7M1a7qhOX4ftA1nwPbC8TS33GrvBVG267uth61awKU8eEyqsZU
AEPAJ0xh8wqeI/+O2IUeFnFi3PQz30Lha7Auae06BaQldPp4PnncAnZP1It8GE8a
WuA3PLxApLe9aH8NjHURQ7mDZnxnnbB4XUCH7G8P/Qyu/1Dt2SOshK06AAbfgvAR
AFNf4JF8XCBzO7l0XIR7hWhc5bik5Yhlx3GeSXk5pv+7u+pAtsaKJa+urwTnFclW
RcvUEdshxL7QGTTHjqGap1y6HTw+3ycl9YFn5PXiGTmWl3gixHX+CLXqn0cFRub5
vyPlLw061pMHl9NH5oFkSWtmkWNZKVi8pdru0U3LnLxCeBUBqbrL2p2y26kIZD+t
579r3SVz6y3kBf2Gpx6MF3W04rMZg/eeZnw6+mnM1dR4KornbFzxiTbMhhcazCdS
KYBi5Ns+glrCOTdKq65MfW7kYKd2/vZCuOrvqc1fIhYS+JpgooufuLDKlZRYdwTo
J1kT/aogOy1xV19LfhFf76zMtXHE6mDdGJvnKOyCJ5yGJJAJ3OdiEVs0Le789DBF
vk2NiSlDcgFIxIAIoMZqXNjd8XzDcuJsLZOgjt6M1MEb87iqAan33ysD2uxqcZs9
PPItR7FBiCurNM8GUyJ+GwcTF67MhhRhJ2vZMwRl4QSf4DLJ44ukuIwmR9SGsXDn
q4LU1gUGF7+T9EYZH2+/up0oYenlpkYklZ1R3m+A9GrYFpz3Ch4ZBl2gNb21YG6k
E2Ix5+58lulg4n/MsBagu/QXE4ln1leeBzxfvP961ssris4AWzchg4FW3ZP/X22g
/Bj0/6TPwoGvIMmT2eM+cDgU2eVD5uuvqtV6DHXlbt7aXi8H6uSUN7pHsBOEJcs9
VBSm20dZgk3OcHv4Qj2jkTX09hOqrsoNkfLdoXV6QLV5WreOxK8dNrfDL2xuVtEV
XFSNvDeSJMk+n8TeWGFqwMfBOUazia8nodetIIPIuojqQ4NBEWn25YiARLX/ksK6
Yf5tmWj8Y7lbdZLu5MHY2rYTbtTswVgZMX5oJoRR2UZ+wzs4BoaHz6LFaihnDLUZ
BovWRsN7QVxh3QncweFJZTJ9YzPzJ4xOSSWfg94S8DeADlqAn9cxw6Z63R4U30tR
3nJ0Jc2EyaxRpEZ+T+gGdC6gafuor6kP3DqLY0IPwuOrBo78H4WwemSH0yiB5t0x
b5HHXS29oG2yMK94KpOh1W8m7oN3pX9HMl4eV5u4oOPCb19R1hvDxz8YPs3gDHcn
tEya7qm18sUUp+tq0MRPwHpuiR9DeSj4iRYZ0XH0rAGuy2pR/KifsxKDPl29QMY6
pKCZLsVPofw3ciKGYDXH79jhHB3iv+NuhZuzKsHp+Ls0pLzym5RikFujNLaVoboP
m3XlWxCARQQWsYWMl/tggLnRdquR+p7VB19oqP15tzDuAIrvou/7qXGvv39za8qx
TSibG5UmNPcpfOXsumFjgoDzAz/oeif+0ODyDlpISWxLwT3FDfYkTe1Bvo5vdXRx
Jt6n5aMxCM0OL+6I/yxWb9V/cEIRikruKSZqlKAAuRNj24NgPt79DvjB18cQnvec
Oc1uL0Qm/8h3yBPx1pd/jqH1dYKIq3Hf1JXSxYdRfLIXXMUAx9MgJuPGMU5lB2Vc
61RpZF/EVGKGJj2B9MydD3oVZZHTOq/z0dJNaU34dgFeFroRvugJnNRQ5DQPQJqs
Bw55sMZdwjzIr/HgYMNqhXzdJg56t9tNZQEc+gl8dKwYqsjyua4IViPcsFH35+/c
Efk+HbVKxyABZmvdHQc/5F8CYZAbj08tG9fm8C0o5CReqXw51hde7Qx6rayQsY7v
Vhir+qPVbjaHclmAyz6dgjEko5igmhMyGahVjQcKW0ymm5fJ0DTBYMNRdUTDETOw
2VPhoJYQHV+V2b8F1TvhnGH34nwLZept1wHHtJglddPyuQRjXiHe8VoUjCS/VaA4
Kr+ETFSVh4+Rxd8smOhtK8n7IW+S07iLPqsPmnlRmXTbRxoKwjwEuEtsfTFIMUzq
BEyESNlDBQgkqDWNo8NuwcltLOvtfDV9v/5ZS+Pq0CfUoWA6jP90eprx44OpSHiX
pG7T+FXtr5faHcWRJMC9rwerfCLNWCRhmzAwozY90tiabbIw4WtvLH4P9/05/Pl3
KUAe1BFjt1AoK0Fr47Bw2L5sRQttyZubaNmHOyVI1brCajEBsdzeUNxAzHnsIzRM
3EupI9/XisJQolgZ7b7+0IzbWVdWDzp6OH9cJRgF9ahfd82gP/09QIonV6eFsUoC
/vfSK2434YRpWhsueMrAQxN7DuUwFJAtMvDms2k1LiG4P70IHMJrBViy54WHm/8d
Nso1KB3yq77kenK2VNtWkVSF4SWzGGd/HCLBu0Ru/t18owC+tzVUO0ePLmvKk9tS
zAYWHlbF0/0pkBT6GJAjcwr9Gke2XeHX1HWoH7e5oiARQECsDab+zc4EUgMASlUJ
yfRwIFVWK9XKuknG8A49UZa/wd0jRobepeBq+vLpDhb/P5YQZ0j4Q/C+ggk6HRIv
7MnFo6wp/G5Jm2soayl1n7ntvnJNSiDHbqQGlhbYQ1Wzh0NM08CifalqslrRbiVa
qnpVKrnOYkPzYF/Thmjbg6pA/RE32UOLlXiX/kfzya/XHKxcQDM4gaS9SVk4G0I+
3CkS2/0uDMBPq0DCcKwZ7SsP7TD5SRCF76z8a6XjMOZqpZPTJIsmp8uGDX9VGeen
9RJnspS8N3pkeihsTfzI0oWOkhYBxvWlwqvnY8+DPpyb/e39DHGSpcp2EnXbTSzQ
TD1Gtsze4/USVATa08NqIXo/SMdvA1IxOZlMkClf/8Yd8tWCZ3eM7QQT3ChEahDA
WfWTVU1DkdLT8wCsKH/2N2OPXvbOltb0PecQUut5AYHcFZDhep/bbYQyj+hKnHgd
4dQqGOvcLNkdSIyQ3ZwDJz3ev+Tss361IyOafgD0KwTVkICxjQZA407/rfcN/jTU
r7QsNoEdDbIVw90JE3KzwbiJqYj+8ZKCjl7iHikyFvchmvVUCam2hOVqY/xdjp5y
UIW6BmuT6bANlS5+rNHhD4ownvOAFcP10/Ew+XFJ8NnKdZ1KxI2vW+fdmI6SOGAC
tWGXqd18GUwRIJpHJ3V4InEmRVE1e68PUxOE+NfI8D/aRZlcjAaBIJOoKwOqnasg
XcNiUpHs7xqZrJnryr4utcw7LJEEWICYdKhK0Y0/5vmxPvrEGAhqifyBLnkV7KB+
GYYHPR+/X7pkUU7wF58FIJ9uiWBIUNYLH1U/Hv4z5q8fnMZbqrroETRtM5Wa5WTD
wa79IjRsa6tYeVjV/d6bZSNCcoXVPJ5jskTYBrNMeO4vLzGftJcQQ5jOILLtj4jQ
VAjkWoPhhVlQ/mQt+jMy3VJvFIe5+RW/7SXFf5d1Zr729oEV8F1R/Hb2xkmYXJu+
JhEY3JDUqzimLzLC0vZIc0XHis39K1MbGbhpzkYl3Oy4jMSv6PdaJ7zAdFAZi/NX
PqQ+0oWmT5RhQb85I5wVhzFvff+cbitKxT21dfMDAtWaWoFmsPSp+0mog5/pwDHu
bZZ1ds962NPxIOjzpO1fm2Dr6uu8YmpIi6cNwhDmRd4p6sY452k/8FBX7s3yXTZi
C4p8x+4bY265XctVTpJH3rN89GQZaeiFAHySCSBa96r8iu3MHrQhEwmeSYVFUY/h
wvpOOewo5TQw2N3SOjtODiHc5Uvxww6Tysv4B08gG/EqCwuuAcwPKABl50wsjT+E
gqRukiMe/xuuKZxKOG7j2dTfhhSjMB6FVRQ22fYV5sJNBT/H8HKeya58H4z4xgUg
KCnVDbCc+3yf++MgmX9Bg2HEcvRNCReNYQ5nK+Uo85U6VaXDAeAnLVOHonHm/SVO
DCidMeyV0l7npVDq/kvgJNoMEPxv73x66xOpl3DpYWnWGRapukN0nmKIWUiWpNlU
Rmxs0lNDmzu9SrWwEPRnS5lHbADdrrvUsO1KXDw0rVx5sGaySV3W/0BxHPZQ/OK5
HKsrE7oTWmboTk9sJWMtPk7KRwouDYnPPOZbS0yW05+fsyRuS1sVQJyIcB6Gsmtc
RLn2ggtI0A5/0qNp91xuErxemNAVai2EG4O5pvQjBrwjECXgSeymHc9EUxue+wge
BiuLFJhOv6+pk5me8P+niZxJRUYARrjxY8MzGIz1AQ9mfBT4IE5rmYJAbIvDKTxV
I4MIUWaAuUjP/k7v/UpizdgEHPWstA/2u+NA8+oyGcf5NJ2eQUgKwjNNQdhC2Z/l
eWyBlWdDUVcq7RYotUIi2G4BiIgqbckkZ9J37RDw/zb0whDPQ73aV2VLSqgvCqCE
QGZmWiu70oqL0IHV2jmGo4helxuPD/2F7ehP5CriJ4XH23O6q9WHwpr1+mFPsCNm
cBUWWrPoYFtP/aLu5iwFMDytHVK9DFPaMRTnKLmYyVeeCt/470urJi6OJMEuGItG
Sx9nL5VsuQQltpm2CrBbK0NyaKXQw750B6gCOlNG3FFhSZj9+ohKXVWoBK3a2niG
rapvgHC5UmfFDPvDKIG0GVm8mnYprhuQ2mCdx9zZohQaOhc37LVAG+sURfRsSEr6
fWpmn50/EObIGoW3bTV9EirTCWQJaGljjvXjR884QsvTZdgm7fKuoTGsyXO17UU6
gaa2TWdP6GXH3bsUysRu/hRQaLxat+LstzxBcQHXt+l6ED5KgpWp/7MYeLG/I05I
txo0Z8fV50quFsjN7SjRH97l8txm8nYH0vyvm1Ipu5PAJW/NbExZ//R6ZTubHe4x
d1Mhk5JrXpra2mZUpCZ9a8SVY8IJgvoc3xsHMYddE88MT/NEZtqQ4+4uFchHubdt
kLpgnTZuy36cJTc375fGzL9LhN4jF8PjRkD2PmAEtTuF0jKslgSaIZCMt4lNPLM7
UNYPSSSs6it5m3MQOrOCk1oHljxfpQoTvtuvBxYz1DIUewZVkBy58A94Cf8HjnoI
MCLDstlncSRI2/bBr3oR7/ja7iC/540VqfRQwQ70sPixTHZVz44lODZ4/mOFiFd4
TJj48r6NghGt4AkG/VqoMv6SLJMc9BeAvy5w5eKU8MSRDTYPIhnuiya64VRFK4W1
VcQVHqUKYKwMEG81A4OI5KeW/N6eOHa5IteN0z9ofHTIMhNukj/aW83+eKTxLplE
Zcpvg89T1Vdl4inLh8aSt87ElxmFoomwMYMe4L3VF+gGUhvwKSaBpbiwUnkHi/Dx
mfzGP6WUanu2zkh3wVWG057s3C80WyX/YUnEGTnCdG+E6c9Z9h7a2fodcGZLgeeM
XdSGmXFQ6e6JN9ae2mAzOD/5tzhq+tCm//1HyzY9jtc2JbC4fbL403D40OsgLFy6
7xXtUuCGXAlRP9loSfA3OxGFS3Ix7eOiV1E934wi1y5c8kdFzk4IzmCf1vSzAxYp
YUfO/ANiOFzj/D/QOKzcpuh2jXvZifxhcAamMap+u1BMUqtAO04n4z+0jqmtFpMC
3xEgx+wCL6N+4pZWPRffgm/5KECM5bTt4Q2VZHY2Tf+uGhdPaE0T0kE9sicLsM1J
b9JlyLiv366RT5RfhjE2mFtnuMViF1xpxrc0FXZhpKTZ4vj7n0+7oLRTZVVLv3d0
taZTllOhddnsh2HoPuoDJ36rAz7lu7/2ew4q7Yw4Nj5aeq/2Weq630YcG9vZtcex
JnPQPElODUzFUxkij/hjgv/rayx9Q0h8ABrHYLKJQaw1E647ArO3g97RsSDnO8OS
CGz6rKYkF08ekw8vzk6otXEGd5j2Hv2STaXqks7oRiF4M7wrXIMv3cMcF4S/ZRPI
1IbtsLu3qzQM38jbSsaquLD/N3A8lLNRMhwz/NxatcTBm+trWpohhkoLiDo9QJTC
4A0yIbZyntgtgLekQ4rEkiavHendHt5/MmKG4Ft9wO31lqYP4ypm1uDNHXoAnIJs
nlb8BTYKoCgqRdGwcPrewPdV0wWBB3tdBCD92hgRiIv9q7YKBjzIyWtj+ev2gxzm
Cp1G/FqJN3nPGfWAd3OHK0AqOm3LpAOSZh9OJtY4d1t0559E4n55v6IPHERp3qLk
HZxtSTyaHkQdHc6UW5a3aEYUkjsS5B9hKZJM/rjGAAm0ec4qV0ullpkb2QHkRY+b
Ma4n1tdsQArcBITJqtCYXdEqOl2N92Rp/x95MbKzrQhdRk5z4J6k1Nm6LKz27eV5
8nzddA6Plfe7MFyzRUBMl3oICAlBAx8D2BA/h+Ffwbv8qo8kRnnVI38mzC/EQzhr
ZxZuEAn+Yq0+wQ9SDTGKeypTwC8301BCuWAxkbXifGKHMXNbZEBmArvejhSjTBDA
TP24RnAUltUgqCZv8KAnxIJhs+NtkUwf0jk3kEBxBSlKKMSy6aZdPD4n8HvJHqTU
FHCqxuFgTP1eefOaGcQmvQ8Jr3hTH8yxniNVGPo1ELLpkTMkE8yLHjyewDcHm1rr
wT4r3XJXu+Jfqgv3Dwzx5dTJKpPEzpyVnkSLUK/12nsjqstxZHjBcqH7gIbvjbCT
uYWhNuRJ5pHhu1FeDbOLzQUNM2w9cDdXgpBW9ZrQZuS6TKGrjIXmA1up2tM7qS7i
IdQfjDkcH+rDO5F7oEUoxP+Wl18Ob//3CtXY/Y9BYLAQO9q/XWuUpLZAsbyhNlsO
FYcf5YrrI9ss25oAK7RQ1rHOIKtjKyGPAV0lRVuNEpj4YiQwKOoOJ8LxQmSuhUTr
wNQ2DDm2DRAnTiXzJ4tTzuozaYlLOfq0yuGP9Lh9HxmmXcB+NMw2KKxmL7W+LS/Q
wJK2u3QeuLAWQCtuPAHGKjQU8XJOrxT2+7ihqtnxJwQQ/QcmTYyK5/Hc9LYiGHOy
t7+3a58cQ/o0gqwiymTctoKbg3wru9ezhwwI7geTltfTIKaTZYyTBf7aa5Rvob/1
tHF5/gJWPvjeT60jteGjaIz+esRofybfytEEkI5GJkrDRWiIzOxLxdzV7U3Cyru2
J3Ri6YULUNVy4cW0/Apk4DKxqs4dawJ0YBJIMzPd3By3ADJArBZUp/tj34uoWRGi
3E3HMVe3BSK1XvoZSFh5eGzx40cb9RSUthkvAISdvxE8j5RzCezQNCT6jQRWK6st
KjR6EZpJqDagUyLFy6KAUjz12QZQDcuMxVc0KUHJf8RB8Zk0m1n0KjsP2Pr9ceqU
gzVDejebiox+mkVb6QlBS2sZ2BCwg2rGcOZeTr398crIbjiAnrcEODVi+succ87K
UrY8gApAz1pKCuZ9aAdKdFBvsfUz5hyBxWoJAFo2qe0QNJ0d4Nj+2PSevepwRYqQ
lJi65NmMpBil+QJcjO1Cr4tkbcyyp7z9CwOEteJgtwnyNG/Du2uJqpluJWgMhSjo
P/lADWn96bYsUE4xZ8PubtkXLWp5Mp5KWtwrFJuU+5+MhZ1tmUSMHmSRIgDEM1g7
kHwyAv+58RiJUoZqty1QGUmavabSNUViXLe1D1LWHrdKPneV1iG3rniQFfKfsax3
2cz6GE46sUdVie+z/h+KDdsftj4dMFLJbYr6SKNLWo7E0VzTr9/hncqrCJDnZkwl
+YS+g2oADyRR3HdPZcRzlmlKaJP8Y+VIqRvddOJw080CBAn9yWJpiyAoF3BbwTI6
BWGmm7IxoDKnZM8Piy9eNI6X9Qh+HBaI2m4YawdGAp3nOlhwkO/r/HssTAuWHIPw
UjM0EK+wXAQyniRRSR66SEJKwOFPMpTqa3bCnkYWbNid62KZq2JJXQIDRGKMP6BW
YjGkndRTEO9gN4wi/GsBfxbPcuUNGfC8c9h9atyEdmnIT2x4hGOJzGz/8CdRbkgP
z3UOtCxDv/lG7NkUNPdB6rPuofnNCeFmAo3eGOi2881MU9tPkgTsofpU5tW4hFmm
oDtHvfA4p2yhmF8Npo0nIdL/JGSZEjpwXR6iyZad9TELBhcLmMSnlSxeXyY9q4La
GX6BljD8VM1ODaN9R3Z3EVTuGaun7YsQYmCVwbvaaCwnZXSihSyyxxbSoM0Emwhb
uXxMPD3l5RKyz0ue0A/v12BBO3nKgg0DbLJu5Tt4M8S3mF/RsdLnhWOstTQ+GLCb
B6YUJJKTAxO46IiVY/dQz940BHJrU759yE4BjQ5cQZFZVJDPQvMty+Rezj4iPxvM
+GzB+hljARsdb0KmS082Ikl+2bqlGAO8q28A12ZGYfNCb/zQTpjx9FvZY8rcHu5p
eGM0Mh4pspc/hyvB+rGDa4vntDMgd5NitfWGqQ078GFFWRYFdzocvidByi78AnEt
6UwZkcexB4oJvEcJDuiV7ngmdvw4KJ1uOIOS9866gRqO7RxPbkJjAF3SWl4/g5eB
DbLreu3IGueOJWPEmxrmueAIo8O78Sw4xswGuUjldtohq2ZjlVyztB6F59LQlazR
JaTSNKjv1EYEaLSC1ELq4uCKpkJcbtXvUzltmqAvIZYC5obdPmPKBHQrl1DIXXpD
z5ZvwwMSoKKhbwmFxXq1X8zir9jzAjGsoaHydlQtLo6QxUofLqG0ixQTIra0j4ur
I7KK4t9icn9+0oWoZjo41/cPwNpd7DSZwcowE+ndfOullirZ4y0FpA2R03x9ZGEO
bLKW8dt8355Bt/nKTxh3oOZcJG5HpqRcJCL1Yu8ybKf+l4GZ2c0TDZt/E+DRqK/s
Z2FRA5wlgbrdnVW9OTiDhXrxep5JCzau1m3BDerWcuA2mVKc2eAyiVU+YdPvsqOy
wWx42mBqBUhEDL26hyh/Q4ZcerbK2Bh+dkqJ6J8RBKCb05lfoJzekb+SZi8BhGHq
tWlHUGQH8+7l4Y2rE5m0clW0n7rKGnOh4/ZddhhvlihQCTCUsrC/27VXo/UK/g3k
Lfu/46i0wCtMyLOLHH1yEMAPkWguZxhf87WhRIXOwWqQME1WatpX/+rU3jMkVbUY
S9GmHJGxRpGHSZuBGQXTlSrunWMpYCKsoJW0qIdLgiU9FPUK3bfaInQnK8g8Mq8u
wnINjVCHvMJqRv1ma9Hy+o7Md0dJwktEZFVzzF98cj3BnoWcGx96nh+tvr0L6EIA
RFpzEmhinY6MpSSBHOs4g/ffaWYQlHIL9YmkPxCtZ5vgR5nFmjwUOOCWiLv/hFDa
zQDSie2lMgB/gK2EleUhFISVDFovqNPYqM4QzxVH7lR6+fPnWywGe7g79pBrekm6
3Prvdl+UiWmXpAfLD1rFAdfbMDRC6pFRY+LpBRDhmjNzRMfZ2y8SZiLCIj0XNull
eadqEu7oEyroEUP8VbFvXqniEblpY/OUCIPLvFqDY9ONWgu+LuixDrZ8xG1WNwHL
ne/QdkIGxcBlevwGjHRK16X8WiWdIEeyJgkHq8d7E2rUN6zAxw+bh/E7J2AsbTKZ
n50iL8m1hwGqVeWZNzus8tAVpuJXTMgsMEQhKvq85G9pobqczj3eHeTnDNBx4ncQ
G2SpgS5fgdPOEFay+1EV9ok6txEQYEz68fp+lu6K+0vMnxE+DvVjPNe1TKr8EWgq
cNLQqg86n4LiF1G3tP/Z4+rZZ0/Qrsuqa9T0IPi9bATHYr6GHeWG1lZizidOLE+U
a6OxCRu9k7mhtgHSPLT7u0FQ+fjZjrBM8NycjadnT2NAoUsl3f4xBWuwLVFtWQRc
uenht+wUd2E3ygXY/y6e4uGec+BR0oTuBFsjbJvoodFdAth3DlLoewQTYONfIZX1
6yDcaI03RA3MeAzzGshty2ixgykz9jZIT7T8NqsrwBWYLehuh0qEEd2BSXqQSbd3
uQIO1HSKmNqA4ba6pXDc+ZOIUzYyrTBW/6NRzqLvsu1uT1pCwtxQTP6Ay88EfbAa
83njtLrUXRppHB05DSB+gizTmcdhXQJBQyXpIVBnWVcA+x6FITeA/FbCXrQ0GK0r
7iiZm2ZMTypneyOQUQTQTvg3FdSeBXH+Am5+9df+ju/NQpqAaN5BvK1DjSQsPvyq
d04h3Oki6BTSvH5ZWx5TyvGGT+1sf17wESq5F0wu5jxUOV4yqEFBkDy9rZBeNY8/
4BZzhZvh+O4kMmr47SMootFQFRsjULIfBhFWETLlTHEFx447Jkhxc4Ydy9BtfTVA
PqQ5TlZnWUm5NuXc4TibyqeNVdQpviHjAo5hprb0zcnZ3CF8se/3dup7i5EVAxab
/Z66jYOYvEJxZ9NmLKuu+RuHewz6GKAvZqA2gRqUy+JM+i1LRXosZfRzsegs4tl1
FnGyeeK4iPyGjY0m6RX/1OmctwXhwduECFemPWKsE60ZvxvKHO34FiMBKjFla7Jh
QS5gkBVOiyFFZIZPGsLgHmms6ILDwpiO+BlCnITOCyso0AbxFXKnJpEh55bfyyz8
ME/Hl/RGDHA7AWkbVYLgYZAHibSHEYIhV/qBfN9Hi9vpJPvjIcZIJv1ba0W1nDjU
oJpcv0xGU4fiYPi7u4QiMX7V9ovBawztU/paTurWZAh5PQZDkbD4r3sXQgecJOeE
1F7uU00dG6gDZ2V8BaA65zT4B+/x1z7K0KnZfiD3eKKdv0zniHGb1/7+Jif+KsCQ
b/22ec7yg3ggTxSDPef7dtf27RKMj1lgovqDsSSjq4Hlfb3muJDZNkhPauaOBPtd
prDmmK3PII2Epv1eSce2teXMlszFwm5C6n/BgwNDgpA3OdFcy1LaDIpw3nFuego+
hKyq169KMDL0RfoC5A1A4RxTZAl1lWOdskH7g/ShW8onkWI4RlUKq/3d+V0F5rI6
IfSG0Y24TwFSdIIpPyzV9dnv1MgqI/Vhf89qi1XHKkTTSxC6C4ZBKuCvQSf54Phn
UoPtEly3KdksNJBnhQq8mBSrvhBC6GPirlMPoVvPAgcD/sZUn5ofcCRrqr7RUa/v
cjm/8CRlt/en9zq76gktVr1zweF11S3vqjkW1d2OQpZZMPihSlQFUDTf2lGi5PyA
y6MLM67RB7LUXqW/ML5oPsFd/SvaM7N8Kt3dNcaDs+JCYAog9xQEwiFS5y6GuReJ
P4Eos8HnMER+n6TQGrVDgaFSJxu7I4bg1q0ESkhOzrKhc3nDVodKfARVPRQYnrg2
jp4O5/XpagYKUjJYOxZDlA2p0YF2PVtQSSgJa02fUPPUwhhMbvvpJQjn99RW/oue
LAFFpcCoXpcshJCy7kO1XOluWu8ahT77eTFgJnypR5MCT7+uQwGsKiUd7SLqIFer
xDJebsTdBg8fNJvxUAp/4/4yYACDCdLVHF+qfLXr2BfoTCtWwHimF8s6lPRRy6wi
wh1hDmQfSqzo2S/jMxyjvgwS0mYSr/be0suI6cDoeSWFrtTdm8OjiPUIJVLojJTW
jmVf83aJGiioSDQjSGcqXHRYF8bk7Qk0vkl4Z/bslbTNmQ0FyPIUH2T2dLLJMWXO
iKGQCyY4g9wRzihOt2chELIEV1JYCRhBjfAjAZoHWu22zmIO/XxmWuf9nB+mGMe5
mCOjamPAF+gwcWfSHniSPYBhSZwaMp2IX1KNoEluBjPEOU6aDgpUYVX2Q1bajWjt
opZLIhOnFdlFW2Cpr63KAoeKQzcjKnxKNRWLTvpDaPelLK3cJz1Z31AtGflDBSo7
KyQALCjtbetRxum4V+rQq/PRG2bZ8CG+7vVwDZhQxuCDrJbwWS7T89jtODNo12Ar
sKQufUEtnLnGM/kac7bJTANTtvzZQSD5cd9Arkn2n9e4/ySMjzjGQjz1eejisXXV
AYqvo5nEjrHsS8jbpzd2VcXERX4TYRsH3n7k7U9IIesLy5HhcBy7uC2UoFFpkKEj
R1svrsV5tWtfifWIH2Hy1DHAvP7VZorno8rz/HiRsWuj9tq2QXoNdQ3fxLXmUp4N
ETDPS9Wuwzl5BnPe2LjPWUki8kSztsvs7ohz5cugYuyL7zY3qDBvDvRIeOLXcy2h
m1DN/E1EkeTaiiiamnzcWmW53GRdkKTUCh1XbYfHTDA9h+dj5Q4dpFPKnVqMK/Mv
HGCjnzhNaAtkyC6xeRQ+ZTzR09ccKPNjtQUTw3w18xhti/9mWiXVQ8gUa6LFVdL8
SL6Wb5MfCvNJ0suzeubCOF5dvvhdt4klkAlTaUuQcC/NBAoT6wBC0mllMJzjo7VJ
DwEYrv8u1ARmzJfIEpm6Z6TbcafPi1jrJGbIjYO8MbAGtcyBuY8v5NUSq1hgQMwX
/H1qRV5VxAgJIlP4WiLcaz6NrTxKAxvEHG0NraE7X43wuV9qYeIlzU6rGl/+7jgY
qqs3ZuHRA6BEafYk/O1ylyYs5b7+NT9aLhtO00lZ3o620bSsqKS+BHUqfnXqhofO
GkSvFgO4OlozKsBr67/HaP7E7LOcJtmEt/PDedEu+yxRDyOinvvaQ46AR4LGE/gY
Ww2hyBTX15+8LY/wMyu0aeg2P5qCg55kLswkL2eosLfZpqQm1DLr/y1/Up5GxPG5
OExfDQqEgK9LDcpREnD1FJFoUGvWkjV2HnD6mdvHXPnTj2vu8zHJ8wx5eRgpZy+b
j2dMQkfftQREuM9ptBTs67bQ6riAO/QNdGcK3xjlROhee41qt04W0U1B0Vd2x7u3
amTaU4/1ObxspoZxF5lXoOIU+XivAJdKlIlgKLXj5v4eKiF7JXtOIuJ0GVSQ2VS7
r/IVtgtzE3+am7z/hL63Fp6lmTcDQSiXjD/wg4KEBHW18gVhyRQrEkHq2+6zarzK
yaXkALD5X3cX3viIgdE3WmKEtIi2RYwzTzfpDyQf5vJt6edEEijfKUt6nMiLOMYa
ZAqQG6nZ708iYRdNBZuzFs6dsPEXf0dyx5t/0+tZlsQUELIoFaQ0earzGH/co+ni
oeGx1jA8IOozOE38Di6cvykm0C1ethJRFv9wdnDawi53pCvdW4EcQGK9+vCJk9gx
IktatEEEqEhBJ6zJu3qDVGoPfLnysCuHzpdQhV8hrNUzUxNaDPX2/uyxb55kqs27
hSGACQgp2Pq83TU6SzCFbOR6FGxf1birNKTm1WzE21WZRkrKYEMGcaC5bAzVE8tL
rFsSdQdpjMLCyTsJHskW1d7ZnAarBTSTfu6seNRLQe+zuUzTwXleGDOBJnE7Osl5
Le7nG5Ghip7r4CcjPGkbHJhpFrEe0EfXJeRBfuYwBbQWbD/hNtLeCMmw6YHd2Vhd
ZfekMc2WYjWYsoEqmVgPJt2i5X+WUWflwrfO97728rfT/kjAdtqsNMiVKyHrtkZs
C9TmoSVpCy59oLPplsQhWHUpWWjr65eVg7iFcX0SxmMSM5C2I/dAH6wXZg/GiAhp
K5DW6+c+hpektkFGZ25KoWSNKfLWFGu0+cH7c1mAq+72xoglwosjv9baHszOfw02
Q0LPboAvWYOjl2IkqHDHUqoHh38Dx26l/ZwhWaAWYP/3bXzXf2GhKHi9BxArzdu4
A24o70z3/f4VsTlApn1V9U/3qfloSiZXYBN3Rv83sRcFHq6NF2oim6ubHTn6n1kN
R4I4P+80SmdMDuGunMFv/H3xgs7SxyTcFq2tXnwu0ujdhWXQC7ZGXif1sQ4A+q9K
dt3UTGD5Eevn8Jf2JzwQMW03Z4VI+WTgWqlzLCONdGwNl5akauwzg2bWtpyNIM/+
dXbLasi9hlxZfc6f+VLbMz8COhPSpoC6nDUdf/TwJw4ZVNmURO9bj+W6E+RxTRu2
FdBHDID+5ApsskPmot2XoX2QrF9Jtc5bG6J4RkS4Do38p2gRNzhyoGCd4/W1xzGx
l4YjhGS9jbRlqHhdpX8P9auS/TFIGz5HlIjWlKcKhX5JtnkXfafNLzGLEM9fMP79
SpDoh5sT9ImcuYH4HJ4KEEF7LtJZ6yhogKgqxTb7poQ4kPMUCzxtr2sGp1ncNKo0
eTtvqTxdynH848O4PcnGoYnl4m5xNTkPOIa+xRpwc0HAveNkDWvytEo3rgE5dJbo
DexGAV4Pwi2vvssbLRUJm62in0y9Dk25HMILZacwJuCYnrVKYFnHf+E6ZQqY90xN
f/7Jko3PtUZRkgGob3X2O5/mY13V/jMVOPvLFhwNgRotaoqgBfh2Zt/k0NzxGivy
K/saFyL2iY0Wa4YJW6GMbBv8uYdKWShw+ao2XCp64U4kDq6lKdpeW9PJyvCONr4D
pPlOGxyxOyW05ACInWzwmfDQiVlQ2+h/4E3zKxPP26uSJRPjExShaG51MUlEVd65
NhGz0qM2QiUC3hKLI3ybEIXC3dpiAVT60yrBza4WpC60km/zEpL9oT/ABoW8H5hO
xzts/Riod4nLlc+qxxq+4a8wtgpJNWdqOO8OEsflDAsuSi5Eg/dLy2UZrZI3DBHu
J/qM7OzgXq2CJJeOxea8F/AN6yAFBX1MiFUlCryBpcRiei6LuYiSeKN+XsvWszPd
Yi617Q/KRIBkssJSJYI0+4erVwvr+kXB+vfLuqIszA9FwHfqTqDIQiMmtXuAj8Aj
x/xMWPuXlL48a/2TtIcRaI/b/l8DRANszwsqLkhsfWNSEuZ3uJpcNpdnFACRbHam
T0JVOywUVFcIq+rNebvhax5qs/eu2b6tHr/hUSznaCDP9RYD5DurOoRC+wjK+sPB
/47UcTJadql5tFYUEoDiGjxw8jmq9NpM52J5k54Hn6j3xAjh3i8V4JFbks9RW0Ir
8uuUiDVnPanVS0eajCIn1gewCFeLdydskLoJJc+i+0YahcNxJuzHXBhFIIQ6UESJ
+vVf0zPwbhJV202Du4DQcuJaYyGhQiuiD9b4OxtbGl4rTisaCa17Mzc1zbsiwNqH
wQGXALk9udfwiKSFqw6Cj7wl46TynqQFtlMgvfDBBfkyV1LwO2Hz2tSj1ShPGX7+
uBBb8CiMEFo3Q+NKOUl4w2XXcTS1kcLDJtvWCu/KB0hn0KWIGXnLVOcB35nV7yhu
9gCqzj0ybf3/uPOzZSUNS+F3vmE59/39MT9d1/Bhy6fGjph8tTrvcG+kzZHGzHm0
i1xARD9u/H0W62R4Gk1aqpSUy0wvCujVe4otXyERtCyfmz4KsTBKJT2ClXEAFnHG
z92U8LGC6gdfaOFAtnc7a8Sz55CZvS5c3S3pVFgcWTo+Xcels+UFJdKsXvoPL83Q
7eLyaqQa2T5f3I1Jb4wuo9q3VYVhj2RVh610qQRFXuXnI3x+qzBApR5c04blAwty
mT03JjDZIN1EZj1Zj0pYi7B1B8sWZWhsaPIjOw/4B3JedUJlF+WwBujsPtU6RDc0
KOrkX4KWUw4ileJ9aQokbv4TRdW/Jg6KTLEgbvFcrvW3PYdOaVTblen9nOGouayg
VpE5xUvMnuFzaTV6aZbMhsKSzLe6ypqzsP4YCx/OwBNRFFx6UXw87m1zyPhKfAhZ
tZB4Z4DI07xedSz73FLoJVmvY8Bhij9Hw1DgYjswNIjjcSpzeNox23lCTirvVrbm
+97KklAEZYLgjnQiaeemqv0ODIn9p7RQ+YDklEaq7sUtHmobHNevkr/OWM9a/AEM
kae2iez9XGFW/GD5akJeWqVbx0SqOfLj43MA8/Hbb6EUYHaArJ0jAbREeyFK8TW/
TcZwJB6/c3Llcwrxxqv24XngbV4jF8SF6eXZ6QUarNwKwhzvSsIVGXBeosjU6Ie5
eayLu4hKRFbY+KogqoAciDB5QUBI+KQhXW21J6fN6dVD7ZuPxNtkpWUIX+gjEjZO
ySQGF/5kBCx6BFnL+KARRPVzvwDahAGj+ZZIT/SRhS7Iw3YN8P7joMrADzd3lCDz
3G9TXN71ERxtPW4TdCzUsDsHilw0Idup68+SF6DvPih2NMS+EaIAzPhJTJPL7K1U
C4XO1TpmV9DY+WS2yXEJY1a2fzwyFTIPOgn243euwJoPwmrZml7QBCAa5ScGbozz
/+dHc1OdVK0znJ1AkBsy/DGpFsxmSdiA24ZPjSPBkpvuEHwBZqaHeh1GQ0ACx3ZD
U8f0hsJQ9CGLw7k65wshC0gxdTMe63oZOs32teX7ya4gCHocIcG8ZkS4pKO7OBwf
6mrfH4QbX5+aWRoB4ZBixPtfNKY7NXOQC/6+hWzGcnnLvEqMSesJNnnjGZehSqSi
uZP/AouYtRA5u4Doav1NYjsVTIbSJklZvbKsx9G7PoZiFJCZMF5Dz6FgZnPyD7Mw
WiDTnoBEhC2q714gR494YKhMXmXqmsB3KPPYUY115ImKSa4qwsIJ5+rFDgE+05BF
zpHEc8+6MlblZ5/hkR5csmws/5pon/eJQBODf26VGPtz1gbZQpA8MJ8kVJjzqSwX
Ygg9NaYVFaqB65FN1Kk4dYoF2g4tjR3vlvtwVL1Q917sxQ+yOw3USEAQTxRWjc5Q
4DxvFTGhXURVVR+MjjPdMwWzQ/23hpx+j2w3roH51jagtSE/C8JvhZ3Szyc/eA+/
o30HN2X9mXS69QNwkXmkKV3LxXKtXaXh5NSmXU7fj9gWLWzHVFwFWlmbfXJ3/mgT
lCHVIwicMWH030UPs9+CoClP4d0JS2EV5lSe5DPtdQNnSw38jpLFvtsMHuX/QZVK
tyEKLS8vhPAbvIN28HjRBAd0ZAf5BxtJAe4TTsE6OqOO34oLu3QOn/7+6h7umbIB
ge3tz5KG7iSyv0N4hjn5qk9/QE6ld9Q/REeYyxcg0+GAHwuCKOyF2YurWT3M7NxD
qy9dkH8w6p9Tj8gx/15j0pydXNqrjKY0UW81eQOdqFVF10gW4rOdRwhAmB1sVBQz
Airw45lgXCo2bJY0TNOAV10FrXgOvVjCYDvxfjr0qCkAfh2meCH7JZz8QyEJ7W/c
lzRGrzcMnsedqOPfVtbIN+ihimlS7I42oSfa/FwnVH915/+FSE5GvSrTUElqEdjm
GpycfvbgqMeiyOJqjc0QlGbIb/OhRTXqJr35MbHPfojBcpHfjgGhOWW8v6dWj2QX
gbhgBvL8J2/p49ta6Q+bANXpge5SbFqrVUhzSdZqIWKDc+SQo1SI1fXyK12qKglJ
SipiaZQejAVDWgLz5VMVMtWvjnTyXLuTp9g+HmTT/ZiNT9nWHZWcF6SV7/G/p2Mt
cRsPq9cMwvwY990bZSTg6oRfMimJs0XWqGXwIr17AH9b/kd51DB4xQnAQRN4xHYR
tOu2iUdfNFKJHo3h9xUA5B/NOIzDyOatAlmGxFrC45WxACk0AkIjbYwojjBP7aVq
gTQ6yVonSgpYw8Z5k2xF6o6y7X/gDVsj9czVm4BIQssA9As5WyC+Z/pXQYI8y32+
KYIWOMD2wvuxXB1vHFbGS9ZpfP8X4/TcW7FnpTXgedpqeobEnyhVp4SwTXR+Hrc2
dzVOC/t/8c8enN479oIqC7LEDJ90zEPNjOAv03yyxCuNhNVe7hK+VdvezOJ14Vin
i2dtGLQcHZ3P0dO/jYNHqsMupMmEksq/70XfKTPenqG9fvbXT8sNyEfS6rsraIDV
Q5aSzdzY6Y3IeRdGjjPZAINzv9cnY/YYqPXdbDD4ms3FgUkEZhE4dwdO7RZOG8J1
KjLM6T8jQlAXRpRFNZjn6y0eL9XDyYwcZJGogusmxZ9m0dYxjdZNBPi6fGOUj/cp
EeQV4fuzFdt3AAvsIgnbX2dbuJbZAomtc4kPWccjFzSMoiNRck7Qwtz7X0iEaJSB
7fXbj1tvCoFZaNGzklYKdxPyKjPll2VXKYIk+O1Sh/41DugyZoZnDvr/PzQ3ve30
XsSEWy0nGWqMk1lqECGyVbYA6H6AZ2ePaSliJhbdCndP6n7zw483c7GHJkm8ZE/6
r2e8nA8/tHFsdCWpge+AlKWVeWe2EgY1EFQU9C7cAnqYe9NG9+xA7HO6cFAc1XPD
2ACDAqaFmyCC3m9B3+IFVpfqszD7CctiitPDZvjlSvmQhv7Y2lXsWFfpvWtlu9sD
u09N1U8SBcKupkmzH+sJRriU0O3mCkhnP05W4vv4Es1vuxuGCfpHVoICItM4YmfB
sv/81YVmcTqA+mcuHqzzzXvlKwRwdVohD3nzoWJSroN687IGU8BW50pAczlHOOUO
WpLOnxBLqm79zeq0kLo1sdUzyKeHtJxldRo37nC9nbqj2S4yUtJxfR8GnxwiY1A5
hnhH/eecY6UJLzLPfKo5KJcSJq3OgJIacBWZ9KTRLtzMCpnH+JyMIX2YEwSMKj7T
uZldnR5YVZXTsXB5//Sr3uYEjvUIT5/PAuGMVmQouS7aSr2SHDkamWgn/+IORAis
jPojlkyvO+Qw2UO1VhttBbKWpWLXKkGnEmTdr8rLIl1OfstqDRl/4wuWotu3N9N5
D9UtcKaJ8KDMWmdU/ALCCjavKU+dZ9vKMixotwrYdGM7aV43Q8OIZPouWhnLm1OA
Hsbu6XEkriQ3VoxFawr3ouSJoZkWzNmUTWC+/SyTC9+NW0ZaQ5iFY9Ss3RPtxfM1
S/c8CiZN7iljJKCEZWsQV1DsTBdogjEcCTDGnpX38xKIDHOnxWOA46CyBUsqatl1
UUIUm/l7N9B3mSi6JJeD3dAudjijryHqXuNGAXgz9Dy4dq9N/rv8GowoG4jeKyIm
JOcpkqoOY9WJRpfuezEFxuhEgTGB3t4OfQMmhMKb25HSmGOH0AuUCqqUyMnQj4xO
q963s5Ep/QNWlPwQ+iPa1l5PT2c9FaYxLGTJXCsNHkg+aw94EY41kDTvrjzWY49D
mXdT67QO/tWj1zrpACfm4SjGFxQTHHcuQ13veSItzLQPKDfcUG0Was7oxBBKeUH1
tht/SULkScEzBnBOtsAxOiUGp+Sz3mfKPSyxYgNfeKXnmyOoUwU4qXuaccvZEFth
0d9nJrzkMXq5h7YLr/bmtklC18EPzDKHIazOXQHsDjkV8s1El7iomySTixMhO0Hd
1jmx/EiQXK7Zospzy7kG/d731dC48SRKjCx/fxFbtK0fpMSa+ZxBISPAvZG5DHKz
v9J5f7zCPhs3f34Y5uvgy3k//1Q6PDNv0AYAy4dD82VW6q1YrZRaCdK7bsnKkqw4
GBjsaFNyFL6f7nn5gXjrVSKueZukJtAsa6SLcW3DKPKpxZlLgIskEPjs4KYI+6C9
SZwmzWLJZ7oSPhDrS3jTXdCTIH06qGTMmTtjLCv1JcRzj2wLkHTts9M0u4RNhv5h
9B3ObdaQYsecXgkfPzaTmjLx1PFz97cSyN9knCE/drkuVL1DznQ5P9PHHY4zFrUd
UpuPOKtjMr9jElZiFf5tdvOYqH7hLNrqNJGc4sUhS1sIbzagxRaP68GgTzaLHcvS
sCIMBx0j7jXCWr/1RGYzwMlJOyAxeFxuXMhGUL/9Z7WcslJqtEBwYsGp9L0jI01B
hdJkgsuY4i85Od0IDZvf6YWTHcvOfycWqfe+Drz6cl3qfXwapKl8qmnZU24SZtMU
/7VitgMSY79nCMT/5TO/yyXUarnfznA3L0G6zAxVwPRSslFpmNYiZYzx5OIbcYB9
Psoy1caHD1qfqVwgmNWST8Zy2O1Z2rf7uRaEa4RuPf36IrCMvjM67CeWPF01bqgD
fXQHA6CuyJ53/cCXUe2UnU70h6mA8FzY8ffSh5fMoiyNvpVYkIJohPsLqYnHxyCv
tRORulXcVRj/ZXtfgvTtV4IeLJV1iW22GiPLYM7jafVHuVHp5OhZS7JhnOfamoYt
lIoa03vN18ZKy9eB73VL3nIZQZzdpbdB8hfFh17HpjGaMhG9Ky0RKALOvuJ7VeGx
cAxzkNJC+FB9IbVn8fdMgT+1tkAddIh+JBjZMFqYWXbmjZgNPOMCtXSoLMLFjkTf
yjZp/qW5/0TxCUFuTcBpXC0/sMLdMbA6phjZ898uODWbDmawV44a8vI1QYyrsMAV
KV0gsJwTlTuDou4IUQ1YpRh2DnCtpZzHukJ61rmhIf/V6/XEWH9p3M/IcUdMnJca
PKtcDvjrwCPnKlb3hNrb/f4StMY2q+GEig0QG27QH3WmqKJ444G66UhiB17QmPIR
HJ0gksJsbpGR3q/IsRYI4KNY5tOnmrUhGPT35qdHwizrQzMq6xOvSgKs1sBOGUxv
D77Hezyx2fdgRKQdIVAUl6c0Cy2FGEQhm7rCDI0ORlYG0Q67DhZuL+THlvsWmYz6
EcOVefznWJqyoL93s7YoOjeKMIOQfva8sjVOA/2P4pBq6V3jibLuShWOP4lSXl8B
0yPYIPzZrjNjCUSwFliiaF16TwXkGpEs1cVaGJemkAp1ncZctJktJtVOkAWJGgb7
grJl37T3neI656th77w7oaM2bTtvD1SDbSfbhCNUcOnqnbDGEkE8yPh4QSnEXAR9
FLApa1wNAoL+UcVECylS1jKy/Vqr58mAKUSRT2FS3GSFS/yBMDgPlnzyEB7lAmvy
VOOk2StaELdqo6fOr0hlhYGgUA5GajrpEU8+L1DedGsFXhQsbm8I3on2wJ3KfIVN
OUuXiUdMhvd1GntyZWzwJTEvcrMGjZVaxmju+5fDb2GT+b158psqSkkWonY69wML
c+7AehcdUxwybE8aBtGZZj+4Y2Ec0KdnbG8SI3pOn6/NiJnJ7aPX+KwPaEpGUjCm
WN9e2zJZb1XkqjG54hg0auoDvvSIJIVWqjvL3kOCo+6nP7hdX/hJMt/awUjk49Nl
Znq5x897idt2PvRsV0r84ZhLCM6bWGq9JnXADNIGJsXIoVsUArKXU1LkhwEOljC+
zftk5Loj70vpzpRJgJpwzsXjw83/psK+lrGSqopSk0OUYBQPn++A1qb+o8uYkA2w
5PfmhyGf61/cPkk8M9gCnJNKwkT5qaYPJA4sdDsRT0OSbRRUGGFWIt3dytFT+VXX
qNkLE6UdOOWN2bnvRvJdyE6XWLdXFjavXJsq2Y21NkilTu2hLNjPJ7FgNVDbZ1S/
SWMArWzz2+/OxjEtiVQO/BGZaPCqTSPa0ufAYao9Fn7RTazaXnGeEMrhbvxvwM1i
XSFsRwOW8Ve0LOgSrnZZlLNlB6atckaOaGzrw6uSwwRFvkUMbfgBrpraUhW11wjt
zaTFc3aHcdBe6okmL5WCTIvMSqO2p9DgomLb2sgcoVL8Tfpp6VvRj2bb992Hsw11
E1Q+anm7YONqlWS7cCFsdfXjOzem7lUWJ5TlDJItn2YHLZPPgobDfHnQcspRKf0Z
487AdRgsrKXPpuCLDisM8lADwhg8uvVICwA27OPrYIsJSIOlt64/EoGZWFcAgjuS
DXcuquwVCbHAVKn73gm1VGSFm97kATORDxgZR81x7XTKu4yv6fX8wJhx26W95MWV
zzMCbozMUychqedprUD/Pb8YZ6rWANqeJ1Ay0iWujIizLIHmgOj18KvaqOiTnxWa
3bmiP45I+8a9Jm69678ogv8Jh9p/dc1QOjbe5xoV/h0LccQ6ymJiyODPHJZMjSxH
eQMGgh7ONkEnKYOtZIueIMCrVlRiQrD5wejGMjTkEr7trpewREDJQaAYZH2Hr5pL
Zvxk/fNUe0obqvMTXxVXdnE32ZAe5mtlMiSThgvCPu/a/iMS90+j3oa/Vh7dR463
+NzcxqZc4wOiol1p4QbY8+Db5WxOju2KdrY1GWVaunz4vab0U2UXAynl4cu/FsOP
vSS2vEy0XrWea2BN3W4Z/m3CxUWm9s6sJhXP81u25uNzVYMH+3Fcn+iSnxGwD8Bw
98AfvWIiubxmk+4NKnmr/giBvab0XBxErGPxTHFkJd0H2smTdlLQn1wBJHPatZJD
3wyD7TbfDkhYC/Hb3aJ6qLWCBpKJcDmyuKvs7FYyYgOlI479fwVhZz0oW7LR3w4r
iSSUd5KM1UnvcFw1uX/V2fNNUHEhgZidf6YwlR6knSFyir62aLxqkDeAuiMg5Bcj
LdpjhtwwrrtJyZ+Egp8u+tfU8xHzEWlQrIsJVsBth0gsr+6aAqQBtiQhvNEvg/66
yAPchIadsBxilfuwgYhUzhKu/M9UigIwVZbZc2OcBUX7pFLG4ReI2i6xHCpa1Foz
VqrMysFCqqOdGQ1Fob7fiMcKOvW2QN7g7Gp6/tejJltuvHmXHQv4T9tUq/P9YWsX
tIjSXtvAddAD4hdHmQToIOs8O2t1wZcae4HTzj5WdiRbQ+evlZwYs1JqokScGXRx
LRhf/IqWd/S5QTPcMJaKDX72BhraKjkVqmT/e3gJq8ismUBow2GGOUERXgEyHTFx
dcIe45KQk+XBVJlhhnNSnX63nUminuhO4IuI6pVGTJ9Ag4IQXG1AsM+0nhysHPpS
CGiskhK+XSbGCdyUQv8yXPg3ule29URYJYSwBdnTJccAWPacjsmx3DsVqYEtsr4o
WgLxoxCxMEnvNaA/7n/T8JOVSmd4XNZ0U3EZEx8aOSslX+hu4rBsjgItCmlPK0vk
vWV++oWiZGm+yPAK3e+IuNEHey0Z0EGMhNdlRXyIpIRKZPWrRaQqmuo0Fp48xWKi
mavz11cWTAGGCPASDZOn71M1aayaLUSxXLV+vlBn/evTUlTYrVzm6dWictSuB5w7
X7n36I2U5xw1FEAqTVUfZE9o9Qf43l8+MgVWs9JbSbSiXSPbnKwVdokW1wAtC7Gd
eO+TKjhsILEbuIgifLRQKfEtaSLivpZZISqiF61Twszf5zIrffkQfBJVTr4FyyHm
VLRS1VoN8P8SkxOHPJVDYr1kAO6Y58v0F9/QnszOgDewjYaY2jrdwRLxbRJYM6hc
c9CyI3P5qvt7vphcS4wndfAW9pDdz76q0M34nDu73IwXRK7ZjAOPM1sZQ0Bx9pa7
X7IAmQrR9u/lwKqGSJvkdSDp5bOrpBhcBV55xJRhkz2LQ9hhFvy5denD1V+hD0TM
8S0v2UJof31RWgQXg9A2EnCodLRJsrNnokcNJXh9cIYvyVI1UujEI0+thklQ0MuT
gFv0IXTvyD5KI9DxDwG3HMfFj8H4S+sQe7I8H9hDHFs95PuIf7FNWzvtEzTwk6e8
QIOjLLcrKvaXZoaIb8bXfheLjlp3h68rMVEp8Mr7C6j/TWTDrmxokXItE3c9JVIw
Rc5Yw5Ukhbwug2+6Qxs3ltOzMtOPfzkfAg/L6rL/8g6D7Jjf+h1kg+OkSLvY/r76
QmrIj7lI5FHVE4nkAhruqcZFuAKadw2yIAg9ZiHEnW/CVEoVgfgfSXq3HqJ+WH8n
Swh5ojkI9mN1W2KLYWrd78qaJDcIHqWzNiAZv0tvykoKp9Nt+f7FbOH3OlcLYlfE
Xin/aCP/D3HFieTtuSE27RL5gYzQVhVtHN/rc6Osaxs57feMUcTADM0FsyRwjmQY
xX0zzJTbbzb6v8JWLyC1ZMXZYlie9GGZmGaDBdjFGWDuB/jQc1yDoGITBwOgjlMN
os+5/uH2OXnRaJM2OtjSgQD+8SfqKOZ5ehONLRH2d4aKUV1XH9yXIC8Cyt2Ug4Yf
A/ciMPr12wrO/bbQ4NWaVQqiNfn5c8XGrQkA9E8HM6LrOEG3B4eWR5ZJ3v1Iu289
W/OFoXeaqkODlWXPheCMXR0ND0xQI55s5ApdrehrvL3O+sEynhH/hFWfySzzgzMz
rjcK8lfmuDtxSO0almuDs+oGeX7ThAKS96bsxjAJChaT4mVgta7OX5htbayPW3mX
IQI15/ThcnglVo60qudrkS03o723M2/4Vean6n4c+MFfiiHUliVP9pXpQG6HLEbx
8nZAUDw1Py8Wv/njJBGFE/fpft+jbaMEhglIWecYaXX4MiP1SPlm3yMPINECVRql
usTY5GvaV5yeG0EJt0UHbH9taEV6JiaKeTHzOWDp3L9apOOJsl7W3hOfHZhHBQ/l
5PRdOCuzPBsh90oAiJHUxZKUrNTv5g2n42Im13RdhhEd6WK0I+8TAZZN3V6xHO7f
5Marwp9qdgxVhFYb/nAx3RDTTUq61Sf3jAIXKskiH17ChoHH/zIVzjEo49E6FhnG
hgl9N/cXNHMgSKBbqoajv/XqnBAGz097MwZHbo1gXuC14feaT8eTQl8IEbQn/BEd
jHCVlioeU21i9ED1RZu1465OKjneg2eqc+2a8JH670sx/rVQZxo5GvbcxwqWqw7O
U56ETPwhhMY03RwiR1tysT9ieeoZHYvcRu5H52yf7ATfO2Xky5FankClsHky2ha+
NKCDXAQswkdKwCoiWKYg8eJS9SuNKCariVA5lzzfUW9VMCkTNcfu+Bq6ZN4R4AwM
JCfjLD9KTRJkAmRJFjUaYDvBbOctusYEtGAC6zY7Mbxt7UDin9l03zmOT+2a0PIQ
aWQ5fyZ7MaC7/JHvVHQoTNXh1dDgPuDBe+F5C23Yhccf0nW3enaShyLcHW0q9MGg
4MaJpo0PpYuaqPpPni7VMGnz3bhYMh6/wZiVoxaRjnGz9pS0+kXnNp7UNh+flbCJ
V4qoDLwNWjsd/SYnSZyPM3mLW3FSJmRbPI17B8d3nYObtcyzei5Y4LcKV1TZrdsQ
WqvkYttUJatVAWYL4WmrfVkQp5ROpY+xpnSYPvHCzOPo+HWIadhZy1oexvL8aAc7
zUbUmvqZXPdVFgKlB3lvLUGUNuNg2Nq6uktRnK2cCEHMIkTQ10mhT93IunDw9kx+
VD59q3xIbVL7ywwzo2E9xk5oqpADKEuWbCjN3+JOHGxRJXxbVuHPI42EF4R728x0
wW1J3Viu+/EF7GYXAh82hDZCr576AgpsNW9CHUCtneCmqkkulHjkXBaplyTOZqyz
fXArZnOJ7M52odDyz40L1vSC9BAApyWEsi7QBvSlyPznOio6zOlhsZEHcXq3abDT
EfAFl013L03W4ebAiUrGB6IQI+ZPEwxCPjN3iSoPvhX0bKIUq8mXsC+Wvj7Btohi
ko8/vp841ES9GqkxaYm+JT8V5fqGelGZ5WxYLyog+r+82VWzEzDdhGWwxLuLg5i2
3z4QJyUFp1y5PAPqYXFNneYgxH5pxaGVaqVwaVNC1pp6cGRkUCp/gPKSO9ZD4yaw
w59ZMScXmErskq8whOG3SwFTXXvCQKmuFpjHY6NCyW/87y2yj7ZZbvdSckMfXmG9
qMAf4nmYKEmdm+b7FMKdC36n1UbWXEXeoh1EABtwuOK4zIaIQHcNymbB95MVzpuT
RhI3v8e93h1LA1WBH5+xMh3RW4L+qwELKdPYOgzln08P+qi8EqYWSu79QbFFQXc6
u+p8bRRUh7T9sr/DQrirpHQ0gaqToT0uwXali6vvg/iT/0PxecjiHtkyxwoNT+7f
RdcR9LnTfmIMBasZyCdCYKKhcht3gSQUv2W0XSM9kDNd/FlXBCMyacpEkdqFd0Ra
2j/ec8RJ1r8DXw6mgQ0LG81Tkx8Bz+yfp0ir+eimeftO9bNlaBX9Rm/QpJj2DIFc
n7WWqS8CJdsGSJVqLsxUVirDOq4gk7+7iuiHFcnrDe54ZtmwEeNVqthR02NkAWNx
88fZ8tmGc96hn9p5zfwSY0ic5z3fQ/n6ZXZ91NFrQRpzJymvNlWUzLWnpY718QKx
O0oV5QScDJkHRj5I6WUjtnlRD98+NvxuKmKoJUjF038KkiLfQ5KM7EEp1WxlSMzZ
HyhvTvHdLidGBb3yrSG00mfhnP2sXFlXgkHVvLDDvNwNU0GN8IclOVmgSYgmO09X
puVf1BhctW9zBTMviM/QnGsMLn2KbueVbJLrTLxx2U08EA/xAI5sRLFe6X8dAZRF
3Q7mGdVWoCvn3SUw1r8VdlnENAsX2Pi79/iuGbVFZ9v8NGWYU4U8T4vvSoKX6MGd
WKnNhd2Yr5KBljAORO2RzcYq/2sKXStyMYkXqq0ZkhCBL+wD5wK5JzvKOkTRSHMk
CTHMHiumK3Qd6omswxBASL6Kmfd6khlKeewy/8nMXLsEoKMpScK4JICZkuvBMYL1
kjiPIY9Ozc6AmPpvIlAeeltR4NZ8Q6BAlNWOb5Wdcv2oCJyRNL0W+xfcVdsD57I1
U042BDZvIkWN+s986tdvHM6e9DVHJK/djmqnrgXqhSAK8hqS46LDKnlMq5k7RY8p
H+uRZqAAOXbGCcI9HS4IRyEonGtYNXT5Qcgppvr4RWXhmwY4kF3LRFZZ74jwNFbb
LR3NG0bcFVFvGe1RGSt1ZzVLFhsYz5HWoZGXgYuKQ5/Bx00nlcN2dHkIfTS6pGnH
TTaJd043OH9Fm7BPCkrdveD+v0ClVnrZ/o2W2mD2XiTGE/gwcETfvw4Mo3UQYbcz
793VE5GHaWrgQ8oDNQ1WBcMNAeDbFiyeqmzQml1kzSfPpSm6NFtbUQ4kccD7Mxsn
hprPDrogZP/qZKoIkHd6IJC/4WlMl3rMI6wohFkD2YMo5XsiwT7uxvSspl1pj5xR
a4EWbVc+GzRRZlCTVYT7l0hb4+hrKZ5LOUlvwS0ixHgt9y7Zn+zosGqIqfhSTuk0
ZXlRCxKA5lMF2NLVGISwc6nQfVD/Ts+p/NuBI7ayp66BVTmMFzN+VhAKOLyFrs8Q
A8TBgB9lbOFoiW8vyVCpTY4/Nhhs2lEs8PkX+MELG97ZNZ3TyKYMRAve9UqxRl0W
7Il/JfwHzSod5SLoVUNo01D6h0JkZ7dXVgbZhVu0SZgL/ypNf9yd2LGP1Xu2UX4s
amXEcOwpyg3WExPu4C5wDs8BHdxNmizcY2eeorsL1sK1rY4eCKDHH/in1GRQ4UYG
SYCILk1lUd0I1N+0lXkIixbHEn0GmSGxptwhGwiBktwffZbzjx+4hpqdgB3lOF8z
QUpO3OZOC6lcWx703Sk4xfVWWcJCzxlA395Zri7yHXmQoYcIQ7dhX75ykhHTmg+o
u0ZMH1NzvblRG0Dd1KmkGWmWieOP26oJJlLUub5Bb+j+6h6DmeSz1ms6b9AxGhSx
LrQZ6zWJ/gzKAHeGuJp+/14PfpVNqtVdCknQV76BuEcfu71A1F6FHkb+EsIvhJsm
oTfaAzMdCj++Vdm1SNMxVQRidLeBFAiMchoeQnP8QIyjAbtlgKt6Bj4PAVXs7enn
2nvSUAgn0dUeUekHvUve/jeX7k8EyM93FE8h6SjsZnlILAoSF/ivulcyqQm/2Yao
uygyNb0PpH+H+ad68cbV9TaW3raLPXaj/Td4lIKuJmcGUJXNWBkBf/Pqrtfn4Xnw
HFHODbw0+3ZFk1UakqfyXE9h8ZyAbWBH2xokBQzDowGlDhti0gsuOBzBABTTUAWP
TmUO9fm2Xp0AGbWKpQDBRiEu+L6VToLVMkDs79k0VWt/pf1xhdqzey/9Y8u9Xg3n
OoR9ZiCr6jFtwD23iBMWbMZxQIUd7So2PM59P2grHTRKXVRHBFr90uOLlc/jpbNd
/WoHQMq/zDXQxjXpyCHPqEs8irFYZB+6h5yjPiYOhbIT3B28BCDrb+6pJFQqTNp5
9E9sSwgGcyOfKOfsREN8EY0QvJXr79ZUqRig/hpdUghObWs+PBrRwdOy7KG5UUXf
uuxK/JH/0q//ZudNcqbr4/e0rKdEQYrjkRHb2QuQMoSWvYYAxORS6Xs/IOdNP5iz
dtzS3daXsJQJaIEc+ZCwdVy9h9sBU/jngiW8JGiG+689RSw1rJ7YiW3IwAjHkfkw
l4ObA45cxG4KxXJhfxDouo10B6mnyyE2VtGxn0UFsLvlB1Y6RSniNd4i9BT8A4L3
M4s6DE8vuDLKhvWiQatGiKkOwc4w9jGa0JLTBwzbebD3fuNl3TTqt8xKThGeLS21
C8gUy3GwEmag3u+Qx0eRMzSR7IwxdEXxVbw0zyEYyFeuG2XoX9IiosQqg2yOH5ks
2lU6KZatvk4gx3Vp5VR7qg87Ysf8twxntnyitcxHEwvGuVIcaqT+Eovnn/X/TCNn
oe3R2q4t9vpYTZ74GFiYJLy6kfG5lh6k9KeOnDv98eW5/E1oB43S4Yor+dT3Ed7F
XhyKSRDtoXFx8D65EfumvRf/C/gUR+WsjirGX1vzAX+fVQtUoTAd/m/YMYJtePLX
z6ikg8K/hsrcbmgT2SMdrL0T3SIBOqO9yRqG1LDHQlpPRfeyM0b9yQP9IrzLcPJh
YrQSv2pQNsrOTVpIiDA2mw3x0vajuY0Sl0XT5DEsBDgsULsSwTBbD/ldFPKIVyI8
8P9j1r2oZroYUj/AtLsUschWjjRKUA2ZYaMBDmNG+1xR56/5EKyF8ZH05x8/HxSs
vS24jy0X799NZWrMWfEsPkJ/HrMZM+te7qCiEL7bp7LjjUDVRHlZ0w0fAdx/VXTr
lkHFICFTkcIbW3s0ZmFn2KWXwRPcUPai4MJufrEhZ1y1kq+y9kzsWeOoX5IhxNp+
zI9wwkI3ukQ83xskplH0phrq67XW66/pFKu26q4e/aP1VTkNb8I9lYPXcXJHfEWR
xteVStIy6Fj5K/JAs5C1gpFgrKSG/RSTFS4RcAbIcDme1y/W5sIRstBoerLClpf5
vz5abAW1d0tTfu+sazYfUxWA6KW++eCluI0uWH+B80DwgvI6mqN7EVmdn+y649yM
tqpbYfVUhU4L2FS1zVHp1cyxDQksatM1nQImpblOoFwwC3fXKCTah2fmbiewXXWJ
ag41zc8xvDXztnWh1X3h/UJfWNpqVF6ZeAwKDQe8GSnpWBBAGkFD6o7PsLCrQu25
HfhdFuBOXS49r+41GAPJ/0Hrlg6e4JOaGULoNOy5+YUSOXo6r3ZrMysBj0f24Ac2
1RmTj5lliwwQcjP4Uun80zyI9TuiMQ62Oa34ppK23pYSO+bE4mGxFir4iZ+9RrTv
D1bolkDuJR+MDBCzMj3082Xi44tUIPNX8CA0j4hg+Uno7azwC7rwi0gEgkyVYrIN
txOt04wX9TrtQ5eoIbjFm4FnHKAwzZC7x2wC7jawlWfd34UlffFYL/syCMuo0Py6
roB9t3e6nhFr7lMqGyV0f2Wuvuhmcu9RHB0AF/Nd1lfiQW0RPXPDI5CZRvXDbyKy
zfVq3fVnGm/ZhirtzZ74DOgtuld9TZjorKEPsai0VxnVolhft5hVnKKyzLatqTE+
EyWOZOFCSfIyySgJQD8Aa64qdWuTZz+2AYoZDEwsuoIGWCYNglem5OeN/EVHxZjH
/BEmW67Z/4Miokx5hGFsSBl+j3rJ1gx/dIXfYsjx3HWGcwfa7gcQsAvm8Pz5L+QN
YCfV+v+aqZmHCS7E3NTZXeguEXBigzS72iml13y0xdr8QbdyJ1LRP2rTraThJpSs
MKpqdHD5SBIO/Ca4kKvqcfsZHgH+8NdemRrJbfTgkEXRZjmLeFw8VyHUocndzRvX
x5cOYArkhn6/28t3e0QNAf8Eom3Ze9bqF/9DvJqnraoiw08oFz8A9K5Qdjd98KBi
ZBOsTDOdN1DPSmAIID227fvtqsHtB2DB5Vii5/0ALt4gb9wHEW2ZHGchcWIq2+5O
7yWEmU8+ko3TdiNgmwIVkrtPDmbWGFgVDx8q/rdFfkv/xa9V+b9UaJxGydL5QDSl
amrgXdqtGIDtON7PDBEWoaZZtxve2ya8cgF3P5ZaDmjfm1mRwuUTu3Kd+yBVofFH
YuiyEMxygE+WeMpYQeTPmY1cYQpKjxdDq0mrQmCjpv2oK3c8WeiT7KLaiHuSZqpS
TWz1a/ekOlLFWfCiRAUq6gErlx1HYcuDlh5XCVoqB/ut9Wen8Sz6+WJtq+KmQyWZ
Rcpx25VwpuuIVw6N17aF73rRUMyoNPRKgeBxnWVTQN3mCA84/j24achZWkM+Mitm
b0Bf9t3+81kKTyNdGVv+adKf9YmSkTIb4bEbBQ47rDpW6WjXVvQwmbG14N5mxKV2
YQgnv3kHncPTUeoVDuM4Hh5wmFxkeyZ+bnnJduLsNLo5dwTSEUai+UZ4H7pCmrzi
f0zH8zmzSB1c2fFjTbN2JNTXtbJT2iGZ/DPMM46laISmlwT3FTyelQ+z/SVPaHjt
rk2ToZLxzwgbqp/MN28wvJ1VCyw6MjO5AOD0MM3gfAMKs/ZFCEHbXLyhHw1eT58W
W9g/IJR4ALFVwcrXzXAqXD+Zs26lFnRUhXhiLb6d6irM5/yz2RKkfdBXuc2kfeEp
LWxgpl6gupRlGPz4LTjBJKvHpFGM5FTD5OpKU7v+IPSj1pEE6Em1fVaFZcHvPOOQ
cFgHIAp09Nw8OW+2tmHgphvr87T1VECgf9lp14QSKkscRUg6nm4dF9TPyy52v3nQ
iSsIxEY96MTiX1uoscgO/is/Yvmi8g5zWwLFciq1EPosm7AagspkUKY61dTsxuza
ftIOAlQIavPp0+HInDzrX5+SuTp9JtWxMn98K0n+sLxViNkj0APg7sTHyvqnliYU
/10pQQaXltOiOwi+QaqUhDt+i5hL/cMcLhqZD5j+784FgHh2eY3mXpCHLBxgE32I
qSfMxImHG924TnNImt1vHg7bCywbn+v1K1qycW0VE91f+TSM7Fe+AZq7Spx2nMyK
IeWVMCjg+cM6Zg9WKL39wDGL7XyitpsBoBq6xlxkSMU7fI5YQ2x5XtWnLNZyHjWS
+N8ANAN311XpyQ/unCAi7qFz4eBiUwc873UhVR4Ak+A5Wxj450KxsZ5LUUpXqgYl
bIHNbgMfLrI0cNhyf+TqFlVcmLNX8cnUAPkZDU4NsvVUlS8uM838IauLPmlB/dOd
ung6l1+RlkOkHbiBnZ4uT18CnC7Hfwqe17Z7faVsT3rqru+A60ChZ5Fx306RIxWT
1kxgwOyxCfSX8G1p8k6CQDQxpjlhKxzDjcI01SyG4B8xYzNncqRDGao1EILaJzgA
OKVEEu0BKNHCthEzMtfdVybFNeODm/L2PTijMYZkRnP9jPxcPfGbHyNVhZkUbFOz
+M/NHk6Rz2cvB8HDvXyEQkxzy7wP+2l/rAHVwHTjTkIthI/sXyu8bl1sbmjj7KWp
7hgZokLLG2BA89yOM2lpChvDls1e0AKcSkhk/QI+SjdBWOjgyQ8GBn7D8bMfg/By
7uRE6fbPcY7f5NBSUo/Fn5AGIIXfphhZsass5yMne1F/68gcxtbsB3bH39W9YOud
6X2juyItfpp6/71ijeQtoZlywPkqBW/CMJh5GBcuf1noVCkC5rUsXmhNHoqVVjKp
4NPzE34QJhZP+q3pQOe1F2gmaCWWYSDRJwiu+/fwa0KZGZB+48eXteIJCrnn6gUP
EtUVRFBGc4EGMs85uX9KlC8n6AI1uNks4aucV1Y9/j1YCO5z3Rb7cEM/m9uXH2Fy
roQVxhRj7bqVvqJSVRbaPaYpuDh9pN20MOp9lA/vqUuK5yU2NdXMEviKzovhnQE0
E6uAHxS1s+toylFRaOXKa4kNEEAGE49atXRAwjY6FsLA3cMKD06iwUQZX7kLW9w6
UhCAnCJJQlyiRqR22r8l/r3ie9QXRVIRxX7NC5RaJ6hOvE5Um68wPEl1KlBZnAhj
px9bmZdbaKLUGbJHYrgIhIWkO8XkKCUAR0r/yxoHUJ9HHSRvToWPggW9jtxXyFmE
ezB0+4/ZxFBy//ZxBukivrFuVus//HN4auoc29YelJnWcbxCe3EwSZFbzqwYj268
V0T97vVY9uX4oB4loT1ImJrtVmW1a/Hid9iuNOwPZD86TUm87Hvd3QchU2/Jk3h9
FxEw5UU8Ng4p+zgUZXrRhlevkZHTm3R/ZRFW608cfeP6ReBhPhjQAaQcjYGLf5iK
8ny7DAqFWAJZbR8J9iro1bsWJn8JclXgc/4iojTdZXPeNZsAryFG88G+3yeJ88PV
aW2ZLUweDTOzTIKjCaBunKz0dbNZu+OunAn4UONED97n6QMDtFu8x7gG8zDnjACr
Rj45b+eGjKpPVB5DgDHb10gNnJeCAvOx9ob8j2Io4PYzxUb+V2/cgr53o+WCR5Lz
g5RRjlaXOWDygpWWgv2579kLqM78HxdVUyLIZZ8afp5ZXrrYoCYHtU8VZ99GotvY
u6dNyH8EEZhTYzpwHdQyOJ//XNG1kMHyugUmDGYLokThu2oFZyUJuwMMUHwYE9Gn
s2uQCRQzY9fKpmk8O2BhslKYXUOJXxo0FMtGmA+xva8Vujrm6k4Optu0ItVmX0Bn
gVdc1+qSefx1vLnmTja8srIsgYW2VnEmQfdEBL+Oc9yPkRMHM5RzTM7cX5MApnRM
XG77Ke1eaPIBzVWTULvG57YBv5j/sFDzj4traq3vMGIFAOsQRjJxrr2rwMV4j0x5
kgUxvNifFm8tK53v2DgmyLhNIFKXxHe3Z2G+mOOohNJv20qDImUiEAc4g1aayUYy
R/VSGKGUq3KXJdD/x4GKrx+MvCa1AU8rPeE6vM4Sz64YNx4rBV9jQ1NmZplUhzYa
Pe6KNqB75OubfoBXOMlSHRXR0Ayh1zWfGxklhMDi59MfHzlS6lTyv1cHCXcSaqIg
Kbipggs9QgDu2ZfjfPNLr9ms7TZOviON6YnQNgDYcioBtC/kG7TdLy9FZrvLyXZQ
H90Rtj8ktmOVJAgFmMVZmqTjveqIm/gUpUCedWi2nepH9hTHIlcOWpx9PCBs+avw
RivNixmgB6cV0nxnx6UxB+bPDhIWN7r5qo9I9z2ZYlGuCT8empPuuxBLAYfNU6dD
zpzPLFMLmVM7SHHG6TxrFaYBQukAFY2JGms0PXjZ0+6txgVYbBcniiG0dP4xHRS4
fCRtHybOVynu6YUxx5YHabzfQFlsVC5FIM3YH4HHz0+sxy0PzIiEd6e57ExGBe+m
Ui3Um0CC2LJbq7MsCIuEvYNy/9dpRSHg+gvufnXDN9tKzwezKbAGJUqnLjOIyfuB
3YOC6+24aR6CCebx024fo+Ulo3S+0By0gROE98r34m4ytFgpSenuB068ULVb6EMv
+e0wWhykEtOYE+DFfIi6Vc3bWnLzsj2hRmnNm/8PpL3E72Ayp2/4Gj1jUYGQ1oiM
zPgP5vAxnwaJbU+NV5HOM7CJOkhgTK/S9zFzO2L9tRPytBik+kMNBqHvnvgEvOc5
xTPiV2wp5CAigVcOkCIk0aYkhqtyjgyM0q5BF3aEqnGkCUm7E+i6Chk9C1Oo0Xwl
ZwQSSduEpkhLwDNa/m4i6OBM/pIy9BM1iQKNmm4A0sH26mv/m537MG7BMJTWKByi
I3O502As4r44WMUPyA9bHFn/XzGMKDmz3v6+6aYNwmi3rZcssvJI7Sc9SWRQJPKk
btSVW6KWLcQFrIPaBLb2qt9MoWro2egGPETDZwIc0HcAZgpMkQjuTkDt3tIv0qFq
mcqsF/F+ISMCYbhkh7YEt5xT0Rh9CPsNlU63rZSmWPmaHB0gYsG3zpAd1J21gp5B
lqZ92aFAPTJabkXJxlr9Ul680zYX0ItkQAAPHxtA3CcxySw2wW13gWnIRnILSlCp
pgya5/P8mVgy0gNBGuLKh1eY4tVT5/+ediotbBXJnayohu3XUA7mEHoZvtXRADZf
vVdUBtJmLUjxPpbZd7cQWGRgx/wgEEb4MsfJIaD2X2LI5ZxZhnUPjyHjBA257tro
+bzTrY1WNHbyPtjIf6AFlS+ErBxYLEYy49DSJ8K+d6qaTx74BHO+2B0dxdJpUy8v
qnFR9PmM3QT//Eh8lxjdt7bmqGzNHjwAI+QTv1G1O09wPZ4GhnlHo9eJo2XRrnBs
g7MLNFva0v+tza+t4hLB5jkvMg5QSe2R0xBrGZPF31QsjkrkDfui2o00xqpK2zim
PyWF2ruO12T0nNFtWbo12p2KmRxYdP83r+Wj/36ch3kDpQrKgHjshz9HwSmRZySV
30VJZusZAnpQjUmeyl3zrsj0PdU3UluXSC91n5/GE5DjUNfrriRE1EVkgdK/+8ER
n4+v/Up/4mZGTdZBveEvV87rdrdB6oSTV1qj0Y30V8X6qn/997M3kb6MjYG9Gja/
wY5dv8gPZZByVFZvHogJLN1vH00+CZRVtjD2tb1iSR6AWpJH5bHmoUwTNdhlBwXv
Dyq2fyspQEOOXUdz+arf78l2iwB+ditKVQ0liddGeqlAUh2KyBQfVuHP257igMvp
N+Eplq/Hpt24rDmbnETBViaqoj5W+jQwJV6OmCoVGcnFZ+MX7AXVwkd+krv7lGCQ
euozRsV4uX3qSaitZEHYatYjCwwRm+mx6QJqkN7nnDAVOeNAaT1vQBmhWW+2UwJk
S5yTxEMPJ/OJbFw20O+wYkFhmc0SZJ6yvEBY0dxagi6TBZyYNcGCtO992972i+6s
MqPv9Cdvh0lSxgYdP8+DDcsoSnYn09QlqDw9QMOUWCynkVPDR6PQJRSthhfg0Xs8
vOMrr5Rjikkg4GCXph+TU9HRX0JWotR0Ej0A6N02iA4yvvsDCRZAQMMaUDrsogh2
gpnEkcmnRhR4qw4uTUuP88UKH/6htJId8Bv+3NMYeehSPV6GmPIw5ZQ48enOt9AJ
i29aQOIcpYr0jLnD8Q0KB34X4eKSh1sBmuvY2PjdfiNCcae/CrYnrbA2rklFarE5
9tNnu42tunewxtFAhjm75J8c7s08EeZ1CJfXYkBaO+wwWE0yhLn47q7csNvmjC3c
pZ08i5yw55qm9YU60hRRqjF6HRTuw035TOOKZft1BhPpBbPtBOmwUkT552r8oEMi
NTRNrXzphu35xZwG/3JqOBt3mtdvbkqR5ierbEdtpsPbAdvyy/VWcQOUWdtjAYEQ
OTgpDR1rEdwDRjGmYqvNzZyQUUp6g/rwLvURirFX9IoGRAXneDyJmePvaQ84mRoA
LaeH8xmu4fV3o3MWow5ZTjUO0be+zmLES2FLKnpX+Y4gUuyEACeU/SYoBAH/ixJw
YADSCMYFukFvbNV4fI3V8LmETz+Ja/u/pW9RH4dO2OsiWlCP95uv/3I5GHbSY2Jp
DD0Odd1yp9QoYaA1qFbYtRs8jA1GbxD1Gu3ysiFGh8txIEeK/CoXGkTt0YU1tygA
DEYih86xVAfbFd93ne/8Yc6FgSDOnO4bELOq3+6vqqaMsNaxTzs/RIbaphckhhlx
IUKTHYW6e5BuwhAQS1shF7BGcxU6ZY+8d+xntPW9qDw7QEGkUeMwpc/Hc7m3NTKN
X5dFPk64Fzzxey2Rk9eHr/DaSPe8RPw2Ffb6xIN1jrlG0lR2FzFBfLsAg7Fi2qPZ
h2QUc2c1gNIxCMYtaTKHHaT53UBPbAw5PoqvNeTef058bQJ60tnMQ5W7sYva2t6n
3b57ajYtc5REL3I5pLaS/CfX8a1hwuzIfP06ai6gjBdq5sx1hHxXEHvoUF6m5e5h
MsOBCFlwBpwNuTctbU7dGYSv+uQsEgufcm4dvxbU4B0va0H3H4Q8wY89Tx4+tBNl
zwyUIHnGdDiZS28MF3U/eDUzh6Dw+vWuiQC5uTQVrod8LOCZt5WeLfCRBB50vGm8
ly0n4Mh+by4GnFw6WU4R2dogiyBFfNtmYQSBku1B6A6wr8SuM8ZM/XeCrC8jEXI/
Y1U+lgFz4RV90nW1tdwuzyiveZEU6tk3WLnrWRQylfzoTHGgdlX5aZhviHpLxN4u
d9xXET5ZthoksyakwFNOOoe2+BjGtrV4VOiZsIrxLof6qJDNBr40STKldHAgDThJ
tPoZbHxVi6iSARIzCYO9m8isKO9r7oYYWN3GVvR621CXVuRzG4r36kGM9zhUYRlm
9bGjzp45+NUffwG9itadCHR/d7nVNmobJXASLbl8Z/sjwoq5WACLxYxglQrjLg92
UdkUIqtScNq3W3GPVp7JgbL403NT0jwTGxWcNYXgWlFHHoOH4Zrn1KjVzecwt4ys
4sPdgHO+J0yqs7fqvMY+w9fPjYrIrarq9XSbC+8yGlSEzJiw7E1fn/i6X/9rXG9q
dCk4jrrWQT2lQbCJ/cCYGYvpoqTNXDj0jlI6StMl6jqGZn/K/nu8ML6kfHAz1wcn
UF7fXoTjJ9kv33GZcicxU9adcDTOFNy5PWQu0UeaIFgdKKHs6UCUvt60Z2Mplq/W
mFYh41+6xfKtM4DPfxzF2/gXd6Rd4fb9/SZx+CbmeGcJe86u5e1fiSJmD1Svos+i
K1SlGNR9nCYy/EYLgnS+CWzcknbs2tYmnUgczhnsnLE=
`pragma protect end_protected
