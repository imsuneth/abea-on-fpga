// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:52 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DUVmollofeWYzXpzG3/BdkmePGNYVKccZHUhiahLZsgwvTOSyO9ODiMS7xgu7Zuc
vPaDZrILh45mxz5Q1wiWsO2glqUDllOYNTQr4xq1BdM3sxWbTbVKoNlEecvUrmKt
1cqkZ4XEyMqizNJGK6EvfQxEhMYMMN23EqwWblth2L8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14784)
Wu2AkkVGz7izzCHCV2j087GCOaekX9A4bNmhT2Bwlu9yYzE3Hvx9VtcxkC7L0qCo
TSQwWKwhICaA3uF/EHaF+/gfb8qhhS5eGIGY6Uy+Q7rKWb52GJkFoO7PFPI7zzd1
UH+czsamz5U8b3xwrc2XMjQBVaVCVwbJ7ZSZe3xFH+IAjr+jCyjs8xhzf4MGfEV6
ftnwL4rI1b8ldbXELOwfKFVsZ38kZ+te+egpGvM9Cy0Z86tU1MFne3+Pl76H0sjr
PW/Vxid0HjDp6qnwslSqthbFw+Fm6OWe+7gY21JD1WU3XQvBhFFQX9vTVJyfwJWd
26RLCk+oTePG3gK8l3+lt3F8vKK6G1Ls4gUWwaSMaIQzRvSK8rzeH9QijcgqRVCe
JPjLMzr4PYgvh5sBbkN81WvVUJ4IevXwJdmkgKSRXAp4n70g7ROxbhVfAXiJVgGF
es5k3NLFOdnN1EU4lVhaJbJ7D0KF8xEvYaipAyRY5tmtuWm0+yXELmy35/HqDNRA
dn8iaMqpyFRpE4vz8ec1Mp2vKT9bIvFLTCT2DdLc48RVpHNZQfVn9NUIzYTzezlt
WN3yEyxwTrF7WWt2s/q0fvWw3sRTPsHTBnvRghIKqQaq6GG9sjwZ47gRMqYxaerr
67MbQqgk8Ls4hKnMLqRrc7FdD0u6w6D7mg8TYUET2e3L7nFnta0KVOIL4XXIZTVV
607J8s3W1QSYkBvRtkJE7lfg1UmU+e15NrynuWIpa05HroL3yEodwehFLkuKhd1u
nkunJv+WOKNBhE/O4zu5Q9M61tVfGBi3P4S/oZ6zSVz0BR112Sjum34nnrwxQudi
CABXSeZhZPRc9Uc2U87zDIauopgxRqfIPztLas1OtiU0k9nnuoAptndaenwAfo3F
oB6vDjWwY5bTuXci2hl6IcZEBmuWvozqGjAoFMak/Rtbb2dc82PApo6dXu9qM4aU
7IydTGlSwkwiNA55PxCQMvs6pF//b+zmyo8ZwPlmRIrK0I1CxcxZuT2JuFyJROrj
NfYgKd4ne44b7ye8JM3JoHwBfiRpb/DlKx/8/Y5ZowfGM2RSXrPqkjMpD9Fgtb1d
25YW0OwfikC5t9rrno9+wuaU17tbVlslePWTJE8StbGPugOLghCKgFnObjlWoyn2
Zx6Vje25qviAOWqhbt4NBAdtgZfKiKww9ByRRacWJFKrylOe5kmo9Eu0YLJx/ejh
4m5dZw0RGx0QQJ0DTnazldOqHkAA/rBx6l5tmujiQxnf5gliQViPMleJe4XS/CKO
vVmQpUaUThkOKxYj1PtWq2xPPB3JHNfABzVL5lK+cfGRlYpGTPi3fteMLcmUi7jY
lGEW7ZX9VejYUsMOse4t0ENDDX2i8WJrEKrf2TzpaBA+WaAvyCm2T7WK8VRszlaa
cSr8uwpRkAC3fR9zmzgPZ6OwcRqL6/32ByhKEosTAO8geBgShxIdDgO+5qVgXwyT
c/4JA4el9W6vISXrwcWuG4IkVwNsMEnCZGIj4Jcrs4SCOsc200EfqvWnkG1tsAfJ
46P+eBwCJIjChoIFQXCgRX5aoxDi3vnjJ9eEVzFNW+psgVQDXs7O+gZjBlVNlA63
L0TaQjSJSwz9zVIbRHRF5yvn1edY8vGIdkeXSqLIiNlM9Dm3x+KL0Vb5uJ9+PD6F
Ka438z8IYQRFtQS2wkhv1FWYGnfp9sVWg+shNnwVjg6nm+rd3U9QtBusw7r7rn1u
iCPj9xh2oHA6Ng9B1pihiMV7Z00Ea9kPIBec7mpQN1kzFkcaWLUM899tTwVmsPZC
pS78fB13bqTyVuD5UAMhJvGSeUTHamHJo8qMVWau08rsfFZQari7pEjAdg/L3q5X
489DAanEDmdtegmH5ZV8DitYGUa5hwF0rX3IOCqez7VJ1QJ1REwe/aGenBaa+dvt
ogXH0qLHaT9D1ske4sB5j49QPteXEC4NcQWg4x/h1lJGvpcIkk00Dm5LWsmOIzt+
MSmxoSEhWbtA0tNibV3UE+nvynkX8+KaUvzA5lS/vH4CzD+aAmlUDRiagtHys9zA
b8wZo41ZhCV6icxhrrfwiDU41JIlfCcKWkEvnofcP3Jtb1AEN0jXB3WAdT353Mbp
xxJX5sva9H/DFhTTwzhUbg2PRazVcj8UKCv+uU0hfpOI1tlExgTQ4NGENcK0IOT4
W+lVuWo3hwQNI09Wt9q3Q2ca0pdP4RjSlZSBaRtFdcDn0PM3UBuN868DY99jdtyF
Wh+8jjm7o0oXLxoRXdCJVk8GtidqOspikupQFDsnNczfSiyDW8fo2loI3Dh8tGe8
9TsYz4OuGoBCL7QxnWfyHU2P0WX5DdJOSSdemBr5ya/uG/348v+yOvvbiIbDKSyr
u/p/4blVWwBaxXN7yTrh1lZh6CrSQ6p1JhVNf8cPs3HO1QMnJlokIk4BqBWIvzY8
uhncU3AnoqhWyKnub2/L7SFBVOCS3jzK/5cSauGMGSLEZIyzZP3HnUpKP7202DM1
O4yMAixae5JNe/Sad4ltXmNkSoZT7S6N8kkWeBLUzD0pS5UDlcRBSo1VRI85SlQs
S5oMvhXyNFMOFJJqYbL5Z3sgKWYqGg7nz+7qcaz1GfvEEBO5I03Y0d1hgze5D2ls
CWRnJ1fGQ924yStAtLxLjtDaTaPCB4b2aO0nOUr4w3Q/tUkTLdfv4us6J/nCFVDp
6HIyzwEqP0FL/edphCtrt1Fpf/6RvAa6KH2fsZxs5QVwFlJ42cCsvo0drqoahri+
aPRSuBPY+FGmggP8AXclNS65vfboi6r/0pv2P7p+Km7/X1KWmpYW+MjtsfAkX5Zu
H0uUWCmX/GPHXJhyH8pwWU1zyIfQwdoLoQ0bejs33+F/ywwZWzRD857bEk9KvCev
1NoFE9iiH+vI4WguB3xDZ2+Q9CxB7D6abSvacyY7GXXg2H88A/H2t49z7e8NkU0l
Bh9C9TI+CHfSvT5XOSOD6NW5zwlsF6IkXKBMEQr+cN5R21LUj45PXawO2wF6RnT/
6saiLrXK9aFY1vqIZgVQO5mVByyEtFfCufPZCzvaCqRjjXUiQnY6lmjlw15VnI5b
Ikmsz/AJvyLSLAj8nnhz2tJ7nEGrfwPhAmyMUcVrh2/NvytcZq+AfDwquB5oRPbJ
TLWudzt73kEv82JFD/NwQud6Hzk3iCwgY3XNnmx2vbn/Mjy/WK13nAIcw9TK13sq
a7CJpAdRdH0KOmH5SMYAtquss5q2yljpEoDegabr48iLXHmjwkuEuUhmBNaT5aEs
J1cKvqJb2iUthN7j9DgXyXhDIrfbXrLUgvzfnyH4Hza4MjO0E+AUoxsHVEr/nI2p
iu7hCybBhx3sT91dgIQvGu52qSaoWSLdZ8hJ6qtCYK9nXWylvst29FNwmYsf+Sre
uKMlJYLe0cO9l8QeJwIZI+eLfKe+XBqJy1ObYHe3pX4HfpnLWndO64aghmUambCg
pUm1fs+KZ6lK9XkNOlVF9wcAVmbWIn3xWzYgLvRKD5EEGdFOyvTDZSLRLtpXL4Wk
HIliHc5is3XdYKSVYIIN76gcJDPLYmOR2N9e049C07ma7vxgBed2SZ+SCjalfOTt
2NmBQdv02BgoW8GIsmFSmTbhRjJcuBxXRf5J6T710/s9kquS3OkTDVykBo2KcKwQ
3dNHAEneeb1Jlksh1QsUIFBIxtd5c/ptbZV+JP9OTEiup9J9TsIa0/r2Id1TJR1e
2WOyaZqkb5CeQDNVreODU9t+KL9mdK0W7aqnyBJRy4OFedQapl7KP31apWo223k2
C4UTGqqAYAGwhgJ92EhZtPqnftn4ZPGHOz7Y8n5e8LK5CewAtmRZu97PeSIpDQUF
kB1cRPNxhW1mqR5qjws7xAqaQbjRx644wU1B5UB2WSzTh0Ed47UlU1/yjQtGoeQG
drA69DfbMJsIVp4Y2U8OUxffszxPPQzYeqdWYhOePabYc0M0D5oZ17AIwMebRqGj
0cJflhOpQc1TuZqsMxny3EbQ5MutXF8nyg+laW1GTgPYk+A2O7E7aaM3+31hVDZ2
c5lbfozycSpKdiGPUbQBOFHv0Q93Z8028ujvH0t8u5HMM3rtqNuAKi1fdcAe/ul9
8BCNX/r6kTBRYn2NIfdAb+c5TOPv3cAp0Oj3GnvH2FU3PhUR6ntu+1wIXccmV1A3
5dAW33FK91+/6ps1j1vKxsmHQTQVflUGpO6H12KvWwK5L//YB8/OaV+ohKfVyYi/
yG2PR78d9XzqDy1FO5/XoXIN4wMeMBf41qvvY1LhAisl+/zpdSZB25KqCVxqg+Rl
Ofi6rSWLnxrIKHdawI9V5mVYziZ+bxa1yqp8fvcurRTb8CQTcjUWQQCt3HRFff3w
j1eCPtK05UQueT9/OWau+JyaW6teLsWjoVHMNaFsoR36dFqRpSYudR0PbQZXrs/V
szaJMywSbEnw6w2j+o6Mp01hXoiBSTaDj8kDi0PZhjYSTG7Ng+y7YaJPTGEDAqGA
lui/ERHDvAndBz/ReJj17jP5LeNKrmvOKHN7ZsMekGZz6hxFAHdMGY9ExVIXbnCd
GkdEwUnxQ2TIozbdC4Pz8T+1FHMwulwWcA0bJgunFk8kYCNiv9quODNe63MB8R9x
id324aQXrhNmiv6UfKrQhfhPiSfZd15qfhbQNFIONSlH5UUMexubPfuobfxI/HqP
8rd3YFcY4EYxo9sRI7FT1ucnsg2oHqd3p24tS26nEBQf/jLZbT9KD6qMuoYoO7Rf
t1YBetsW27+7U+S8JMccYiJs+CHHbyFpX2K7y/lOPLh2Zi3lwfN0abWrHlzGaFOk
W1W0XfOSr0SdRa5RHxTT1lAqBFXdZgNyeUC60vPhOpjRI8/pOrkLQnjfAXkhE2Ik
ATs0u8K0sKwO4uPBxybA5++l/VGO+pWxGxfhkvJXcyYJtsUJ5GojDrMMWgxklYrn
q0WYZfaMBJU/emLYdq7Z0E8Slqouhn3UQ5Oz0EF39Utjb+vqzcizxPkyea9Yb5Yh
0NTBa623uMxQ5yf56wHq265KknLR06aS25whwK4PTyoq5ERVaBioOk8IrU0qGp2H
v0w9w9E4H7WhmCY+rG0VbXBvNK/1jfSm4OBQ0b9LSA+D7flpUNzXuVJ9kbXYLqjN
F1Pmoh9+EDBOlLq+CWfNrUwYzRvyKdWGCQMjrVvZrBA9QFCTTmpMCE5J79jTuL67
z25oX0cBEBqxc3loHQHrE2Jn8CiHUPjyjK7s0m2xGBWcctOGtxMxRc/8yzPBxffd
ZrEU1R7j8plrugZYGYonFfpextprVFNsDvZwj5FpCafHs5tTfx7QNVuZrN3/b7GW
JJ1+fzpWMhouEjLs9N4VqS8HR5AcjqLFvedO+ng7kg2QTeVUW2pF+zstOxj3xJM+
gHwQsMeACBq/BMhwcHThsbTczBTl/fiuC/8+NcxdtGxNNJydkWtHje743KXEWFW+
IsWx//teBYxz8H96G6HzCCB+y2Q2oYy01J0Oj4iNzUHpcKpQiOj3IGFrbQxeXKGF
YCiCxcHsB1hNx53L452BkzlKMZlDvoZ2QtmUVIXKoE8AXp/vKmXaNzT64S38am0q
iocV4X+exFLLDTRZGybRsUZIMv+yCA9g7vYV745LTGNjfXMPc8jArff7zx1wWvYe
uGOkhUK91xf3ZJpOzOeKlqzpHcg8wDhUjtGwm0ApzwuIXJGNoh3VxzppX0FpOg/g
gDVnHFWmf4gKyBYrD/V7xsKvk+pKGck8XJZSTQeru4wiWRvmzej4xa659LyWfc1B
8xflXo/6SuJy3CcGvGZShbaLIcuc3VTxe19/BV3F1lmeRyt+Me4pQjD5WMR0EMrJ
QOoAFALzKyrG4YWZ0MsYMcAda/QA4288lx3YC63/7V7ZpUGw2g68caQ0LWE/h1/K
7p8YGVB4jLfTsOy/ocpkBCaPykW7GgRSY4ZgHccZwPMoNaAfKetgPjkCl2bLNCsO
yPPLHL28wRs117zcX9wsa2uP38MHmUx4ee7CLjObWwKTB8bPWjFBMwyzlP3uoV/7
XTooGaeNkCp4Jgyv3rDtLzWHve3yIgyJbTZOaq5WlGFM4DCGEgfc0jKqQNSaD2X1
lmZuCxxIx5g5A/AOHA+w9Fy1FJiMmPNjuP6Hm8PHwBihAgzkc82jM8PSKWvIUK1n
XXJTAPdID0krYI6tvrCmMvcgAyBeQfw3Z5PPFx7xLc4K8xgQJi+ycH0I4E7m9ejQ
rSzHUQTKXAmlgugAo/43CbZzv93Pkiu8uD/cCaIrbt4t96GRYEOWBMYnr3C8BoPr
vVAbc8Ltn2IyZA475RLGBC5isv6wdCKARb0BG1Ye//D3RRXVIzmfx5a2pLH7D6iG
TYiFiA7e0GEuNTgM21tsXqUcaw5SNzSQ9wzeH5LfRYIvEGfpSPTbMIq30DCvh8l8
i4hNYrmMxYnJPNxaZ7r/eXf51FzoYs/DyvGvPjrg7g62ZLEHjjPLME7e6I6dzpRT
Rjw9Kgwy+IWor3kHQUB9i9B6LHTrZJLG8fYYY5XeICzCtQXp7vpj5rpPPf4uqf5Q
QX8RYdZI+XDFBLYEQUi1nZwjkq0KejoUFYQnSurXz7EstsoCG7Qr4ZJbtJRzHZVr
hESvr6V43nKmi7N8CELtKQEb6yUYfMvOTIxiOfP9+GIROWVk2WhOfwMUdFSODzc/
VPu+Exc2wqMJzMGIgGBPsjluDvXiTj/EOT9y2MtJSgIsynT7JdGVZniny+JPhr46
QOfYq3nC+TdRc1zBZlG8N7LNvVdSjXnVG+MvD91IgMxvMA0MYtfyLdxumTg+Q0c5
ryKE+iE1f6vA9JqtfoSelmzmwQwmoMnsSVmSJqJqfFYrfASb6GF61VzXP8p88dR8
2HxMzJ3QpURHiEicg3ovJMqiK1wHD6Sheyw20Wkwea4RMAkVZXBq9k4bxBNzCOCU
aUVF0ajKwTECvAfTTrxD1scF5l82gpuyYDbJwvQdAUuFDstUzSMuI1HzTWwQvI7P
j9RWO7Ywap55mCLqz8aNKkeNc9pIWwUtqQFq/3I8SZfU4UtSqgruz9ZGEhH+omir
JpizRxwMUzgFRxj6rYkaztXoio2Hz1Og+EYK4375dpmST8joERJMh8JZfxsb9Kis
wihgwgEHb/r9We+DoSvO/FLcagC617qU1sM7iIUEz7OhkbDYjUICp/GZBE+94Fmv
7LEkA87rxUUlVLiA/cpy3ZsA5uHxD8UVS9uIqLcEIvFmDz67YKy82I6we046uYV9
jzEi6QngNQZRA3K5ocQrP09JYaFSeu1zDLi4PwjWlgOqOzp4yfMaLiB8UH8AxZpG
OXWcqpKD7h7ULIGFQuTNpkEX0453QCoZq8OP0o4aOTGL6npJTN6VnesvhWJ/IKGB
bPOdjsw1pAwOdYSo2rgmY4iP0Oof5zlGTH7Wn53ld7WEST0LeG9SVbeHdVJ0Klgl
wQuVyKhtbWFyjWDbPkFH/TwArcX4pR+ktm4M6qpDbZZj8o9WJnlTbcVh9t/GLjrX
LppwsP9K3nahBsghcUEL/f5mZJx07k5fBFvt3cAviX1OPsiqEljWXCEuapQTbVAu
BC1PDUZtwwcIbIWAkAthAeHdr5+7IAXI5+6Hww/3CuIRPJEvuYRT8K5t+fUBbfXF
ewqBbC2NJsvUUcDUgZbNgh7qRxanEc3lhqZlMIha5jNZoQLxOzoF4YvZaJQhCSIj
YOYuc7kmWHHa9XI8R/TL22jCDegtSYi77R6X+NbEVbvFL2vyhq44eRtyW8HPgP2/
wsGOAKdfSiusQ56ihQ3aBzGuQF6/MzsFM25p/ziMytJjKn1x7IrNKRwghxZA//GO
8pWk687CCjIDesOVZxKDGFrJmmMVrXeATkzb6aSUZigyMWi8saV5r6ibzwKqFn/L
nTSf1CIiWTXWw/0Ri7Q5oEaGYJDMIPcF9CVVnwKiewU7UF24RrjXV/bAknp+ZH0R
vh0/4iQzNePbZFqxr8H2tlKUFLBTjoED4BlzGG6jt1fH3n9PBwPjLS1BirDUqvju
JqSZ/wJTatR2qprKpMZmHUp/eFx56OtkhEeH/1By7c9dPBN3kk6k6LJl/DWYoXfN
2GNtwUVzTJTWQyl89luvD6xURysEYYoe/AuchtN5EmvxEe1zIMzyJaAWa2Za/dUM
te2O3RK59RuFfL0jiKLKQAH+1KML30VRSqCpaGRudEX8mbY7T9lkR1inysw6wzGC
Fcms9m0m5+F4qvJ+s/Q/c39fsdGmacIx+FfIJm5VSPRbYNc5b9RADW17H7nXvIft
Ss5V3MJtjeq9dWAn8vVrQ5l7rKC1iEVLyjZlSRzMzyjXBznypWhCS4Gr611zwXwo
N3Bz/2vGrBBssPnIv4N5PezKGl5PqZSA+6dsltWXC88x3AGj48PbaEpG16nE8GQd
Lv/3KNYZGH3hWJWx/QX2cruBFIgp1wZCc5dZDSHTYhwVji6yiIUh2PL6BPQXXmnC
3/awDOkuGklUj5TTtamosHWFNWS26mXFu026BTdIHcQJeRUVbjGR98VoWoLwxWHP
Sc8vdbl/QlDOp6z1/8Iy7+GzUdz+mQM6aVf2me1iVvNN4dsDOtz8yZzLvrqrwocz
5pqadsyaJSBcdCF9ddvesMVzZks551Bvoyiq2tHu8DM0KARwZbHIyEsu8v4emhrG
QaHSJwm7m3vuzaAVKvDMPQda8uusmBW1S2v2ijg+uBHF0soB5ASbxvwHJwcaDZVZ
iO4GjDFd4hH8L7P1VjOg4ifaT16s8TCnlqpTLO2+G7yej0/O9yTrf6v89J+KFrL1
+B195g82vAiBOEi/fusWUjBUswPW7v80K48q9Cmvf4bUBhSO8VahrjdpICBp6Ttl
kXgnrWjIq8a77ZG7fMJp2FJ8k6VWKvwipiOmaDqFsXvnouVeivhcgg3Ib9+oZgnq
LGv8p3FL2oGr0UDYyP+u+FHVzKm9azotZO3HxveCmIBItPBIu1GxCzpKWHZo7VE0
zvo6zUSjIkMz492QgnnoO0nVZ0kBRQYe87faqFsxdtUQ/ChwfPrOJYfRLqc5KIKf
G2krgPR3nEobsAc4kwA6iYZK19f/ngSJXdHGJxB2wRJmPY6imsvrb0IfOuCW+40l
EnakMLF8guhiIfldeAxwCbU2YKepvMzlyuCFTFYYl8c/s+adoT9q6Yxajrz8a7Gf
HdU8BY20WoU/iItVzvt4dX7dqORWKXOzVkl3P2fe55q5aHDY/o42DToNswHCCkCf
m4lbih2LowZhXnlhV0hxpr11v0VGMTpMf38UGy7KmjBEIyG7vHaCyqpsWARJbs+j
O/lXk5E/TMVEUZdr/7mxdKuXw+jfyBcV/AqrSKydXuEVQA5SIWzSa+tSaj4e+Sx5
lHRMsnHOLJrUj8zjgE5jtBgXgl/RIpwkM5uZQwo9pc6JHEcA0CToeo20y5Zv+GAr
WF3pQpfL3fLjQbt1SKr8/s2Ilq1LuzoGrMHbcPCrdDvl0kmgalTIWGx5vvPXdmc7
qIZKaWlt1EWR78NlvdVBvYJqmRzwGN73jSTxlk6rxJKFF82VmQULI279E4jQ7Kv6
aMftexDc5CpCf9H+XPI/QKTXeZE32zIgnI9ILhvZf3gi3LdKChhP1YCSLb21ciE8
UEUcXgDMQWbKpYrXDcSkmbwwwJn+tBY2Sfr0/d33bPK/nH1EFbYIqXDKHf4aSbdI
XSm9kMT8/AURHSfnnXubjLkzycqcip0Vape0FgSxmOu6ruda9xP3+wCBb6/qUhFz
YEBaeg7WOOWrDlWN/2+KBADSitWjh3wxt7L1LH2PwBdgC2fnIvwOlhPpd4zPbid0
yVEI5Qu6UteWkq4WXcSbFCHJFB+FcNa/jNj/hdDbqfF0xT1/wALFgPsyWjj4pVeQ
zoECm7YnHV4x+6wJjmUJtWX0veL4/36wS/QhMzeO/6G6nZjMMm1rmhnh1EQma5or
7fjeHqTNkO/5/SM+g73495umvtl5RR9guEHdQNdn5wXDLCiK5DZx7XcL9opboVZL
QWRv0AHF0+RLmCTwZ1ec9aVvfq4YN5zCuGJMsMbY1O5bp41M8XZH73IoGMoFBOGk
o7bBx0bWr4IOhnirVNbTGilvAK0wZff8fZHsgpvXIn/GZJjfj6SOaEv/QWV5sKV/
EnVjijqbbE7vy2jAtbXp6AYR3CV1XkDHViw544WEOi71+jctVpzVJPpvGRhaJZJ0
qUInNRT5khfEE2Wr529UoCOLL+Iw8n7LuNcFOFtvillM9X4t2eGMhZJW0y12d3qg
lBKj5VJzu80XoyZNQ2KlCwm9iJJZkq053Q1itpWGvDvLi0YLx3hhmPoSDcpEa+sx
Hs6PShwi6HIKGBlRj2dlun1b21es+AUpnOillPhLC9gCjIiebKenF9TrUJKwBZH9
SV4UZAd5fL6Zy2uarB2+gaFuZoA8o0vdLR941qGWvTEodXKjJrYyKdGlY0fXY3ce
IuUoIJFcmO7o9YQp6dJpBZc+qYRMG6LISTFjVOTSmjoHwGB3IOO8trpk1/kTqMyL
089P7HMZNv8fX2NkbD2v43cSlGFTS7AGYzRe1dVDwkexitubI3rBNpNHcx2hTiJM
uGwF93WA200KfMaqoS2HdW0EP4UvjJ7SUNP3lSqYvFrQ/4Vag/4SZhOB57MfgZx/
tHwRzRISO1TkhZQ5R2YhK4PaliDbgj/9x28VeG9SZAsF/nbHMsHEn+CBdY213XsL
q7WYDxj65Ae4IBW4aYBgWLR2UM93fYrrXZ1zH9cNPzsgvhvEG3KJgIos1bzvL87u
08yaGXLbd9mNud+rPK57SdoakTBwfWwzjbw0/Gjt9A/cUoj7fsAjtJTwkOnmrRYu
2KvZBa0v1WujoGD/OK5Ycfug0qgZZIGbKjxa8Xu4BnWYMr+pQ4RDZil8/+XdAJKz
QIZoszusUIx1WunUU5q6Eflg4BfJYJS6RLkKML8uWPgqs/3sLxmeQJGbeXQrZE17
MyTno445MdKLtHW4vYItMW6MztfV5KHRttBr4t6ZIeRpwweMcfvGEDZXoGfQsQmL
M2ihScSO7UUYKR+z2gDTvNF7XJApOIbxU2F5AyNP+P4HrNpb3PSHDgdL8HdOSOzv
8Rnh7/7FlUq6532rK99OCxaAgzqZ+KlLxCnqdH6Q1czP6armLgIFWvxMlCyUg9Kp
oOsiQm04jmHjwWh1O//QVs89CJbZOIJ5ueJLPvYyUx6PJUjiBw/rf3S4XdB5a/Mk
JniV88TiVZa9NispCja/miRWT53hNj7VLOMWpIE5LAIP9f+JOfpyeBdm4I/7sVl2
83w4YKLiFuBgEd1CAdhO5GUZ+rYfw7sW/6DiC8LyckW5CFa8MIQasR+wBjUEP0D2
GFgaUEnXk+r4HZ5ExxsoIQ3R935R4xaWmpPmFjfLwC4Q454Cb/fX6FFratD9Owv0
AzZuv0KTh2lPU86JBPdSUOe7KJ310aeXIa5G+riK7+C6EB6Kjy1nTN1zPr/txbfa
3d2Ev4CLRxWZkGYMYAJ3eJA8o+ELgLI5mcSguOeGbPZQRsR2xuE5R+3SDAwnBrMV
DTUStl5+iTAZ7ErLRmVvQPniBdM1Osa1Sf61yrwqXJos7y0cERhmrj2ABbquizrN
XFDsNMyXLVDjDFSKn89dgRR5KHnVijC537G3opwJfxvp1ZCMl3KTlvJi+Emk6oUj
vjWEZV2Wl1UM3lbK3SR+apFw6j4nx6u4Ig1iDYWYFDMe/XbPnY0lBamSQ9oh7/IJ
/KxI53MpYd7SSxtVEhDScfe54NSMFalfOA9XGG7MFq1KvblWqypfgPzhdTwZzRCh
HqgZlui8HAs7U8rj+H/kQFSGVRqJBQMRB5fuj6ZB+ISqI+udE2Zs9ZW6T1Ytpd8V
1i0QPPjEJMt/0w9Rjd7fd5K3uCfwjTxUnz26M1GeeCsghkH2MOgiEPtB6CVkuzMB
BT4Vr+7ODIbTh0LQK5uqO7jMYg9T30SGT+V06Ds7cAxTskKIe6db05ltPE7HHlsA
qWPC21TeF4VziOn/LpBSTvdh1muuwYvBLHQfknCMjL0gS+gzpcDn6EAxF9i0AcK/
jPBz/cjzyjY6RLTNhDsmrL/N7w56zazsc++I8I/BSDGi6mXzlb+M3dV7wMf/dLrl
Lo0o4GgJuzv+CF2yFy9o6pz3YrpXFZkf5CaKXzIFadB6CIqlVYTK+EakA/8TIIHP
12TnHpQlxEedSzSz59m3iNn4FHJUIvpvPhCUaY5e6HDLv2kc/WmsaXRJTw5GRiBw
RpfNIBZ9SkmktdpI9A0+tE3KxFTI58XuXnm+zaSIWr4hjABMMGPDWUTQx48OgbCE
ppLr/nce+gZC0ADgwdt4auyezOoK2JVPqc5+rUKkEwqGBCq8rfwBAWVK9Sy1qeLb
lpR0Q6YtMurL2sfuezt1W31BYkUY7XfY3feT/tNWCo/+3b8icPyTSH7Z7o0ll17r
qAhBbdBFD42Mz7vvrQHJu6EwRBEy5zsDICMZwfvCxBMH04YnsjlRo5oIlnCPI2ez
mCvM2JhcbrT+qbUwWVEd1eOWFp/3rPkI0vobdEOhb4WZ8dovLgzVATe6SqDhsl3n
E0HnE6VGEeXUoWh8pEMXSxxNTmSDcP9gSy7tM1RU/ql/LeSc2f3E+NvJV+wLRCo/
Iu6dN2nDeWY5jJ0cPJa9mrERxK4wf1izLY3kPYMrQqNsezTt2Q1NPXdH50ZOvmst
h8lF3i5mE15sv7W38au836tjKWqpQAg+igrPKCl/qXAHrZ9JXuUBDbpNugMprLXc
1HBp7SkE+MVu9w+YwnTYF9W0vxq3hVJIwt/vBPYpVVpdvk9nCcCTtV4uT7XuyN8B
Icqljhp+QBBWC8Na4Gijf1gPvU4EnBK2DucgSeeWhcgFYm4926T/pbLhSXaysQlO
G9UoOunvG4F7oTfGGbTV1dGWNPE2abs0KmKFJHC9jh0yuWB7i9twcJLZGtra81m4
X29jOOcZM+g1ekSc2pVqpyiNcDrS3ehTWkSVjecj43QNV26art7OjUgshMoqa1pj
PebLMyR8IBLVJ29agKhz4aJK/vku556Dl6ulpGBGOAfANHTOpXG+h3p4aHaeBPWC
edoKhb7WLG3hbswX1XyN2dO7pT5L+3bPW2tTMkhIVTEBTRjSr0RLnidm8m/bmrFp
r/kfriwHeMnRyp/9jQ87M4tT+yo285gUtxOujKON28wMmukhM39bAHAfQsxGCOBv
+Bn2G9Rl4/9hN1ckNIMJSs4yNPVYb9MRkBEYmFo/iWK8/tPiB1IrdxW4v1gRCz4R
mvR/bPaKR3gk0TG/Yaf4fw28h+et8kECZiWjQVOdzUoxsT82A8W7o15ZZD4vMdyt
AZBVrvR4PQwzGsmW368Zm6kxAKjtkWibf04YhUVBdTwkBU7AXzhf9eyny5JRrwgi
KkSlDDYJfzJYGfBOYmauGqFBzeganlGTu1IqM6eeEtSmnsTZ20TDXn02d8XDuQs+
T1YVPRBdqvDIhlYqXnQPAjejr5m7j+zI0hOzzP+mWGYr28yzwlC7rhZ0V6z1nFEs
WbwSHyJWqxk0s6OBalKfbyLBPIFdpBX3VG6b0uNNXina30XpG4Gk3+CCqOmHK5/L
0Xfw0UL4SBN7S7G09qLrHBAcll5jTITIWc0WLcBaBv9Jhv6eWjppGkLN7ciW1z6l
8ZtP8mG72wsvjXjBTGYtLCa0LdzIQ2k76SW8A3DoRQ0QDwmv8rgqs6ifvMzsPGZh
o1oCpqkyeAuaF8omvDmR1k3pcgp6jk68BYcAIrIOiOBi8XVtWDa19vQJqXJtvJ29
OOMJEpmtg1dwoMbxTRPzPfjMW0/NIc9n3rBeiVCr6io6E5e08w6EUGo6DdgQC1vw
KfG03mvcGsvFn6CXTtvt5Usy2GETc4R1yeXkSK3x1sKPeLtGY/7C3biwDhiYX7M5
XC0W7EkBJ1b7JxeEKvhykFiwVv4V+ltNZy+hlzgjHq7SO7+2564fVVl+j/+sobWG
l3dHWD6e1pfRptvmLAXa/A9u/naM0H+qIBNQUUaN64DfNGhtd66cmVbB1Tq8N1Tt
DsCOjRkBMNnDKW71jQ3ldlZc/ZrbxzyzSHLFwLMM47PwBB27/lu55fMB8v5jZUjx
zNgKIVM9RlrTBte5bajb0TdK/xe2z3D54FiqwF3gtdD/WJGI7vEoZ6R5o+zpdwJG
BZZWxnjK27LLhdcrRsEvAH+eNDWSJ1pxaKDVKRCxiaV/VTyOAq8lPOtT9lI7Y6tA
aZj6umD5P8qWvHJR/sdu1Seu2UjKVXyWCpbucLKs99TF46oFYyUBN+n2dRrnRVhI
MoYezbmg75veaA+yIbrnLueW9TYdPU4kVL02uYAEExIOcBIlJhJKYsKvzRkNrm1L
iNOcRfFWJdhXpThMUUlU29Fu6vRYpdUGmteaN1U5I8hTSF/gm3ISZB5qEN1m47EZ
t1m0xeaAgg9j6VkoIO2DBHxyc3sA6k9OLFTjOY+sli6GlNdof2El7YO1jB05G+w/
p+LBNZ5P87pNWKgJGyer/8EP0lvTDmomWDQD0HvWTcHHDLXpaNZnpXfm0IbnCecP
0QMaVL9sY44/KzMB56u5TO3xVIGLFPdqVHzjvMkJw210iUOtDkgd/ZSYv4x9hLbf
inoSXI6zRyQI3n8rejixYQiN2d2Nm25B3V3Pc03lR8mIDKHnBzj/DR35oaigqXI2
rIYLtgwJtqe21B1ryjAbzo+whrTjKylz4Sda5V+TojHZBGLp1QUOM873C527IBS/
gneSTIEhatLrLbQL0R1VHLuiTIMk51FPx3XaO+duDkdiO2Xe+Bm5c0rl+r1mtXaS
7aEnYvH/uh0mITlb5NK9HwJ7uRS4uKT9/427bJlZmxwjyHUYfxcAWbjXwqYaisKD
3DtN0RRhX2FaXQgt/okm4W5Mdib/JVqovCHQFb1fHbP5ybULl+RrWK/nqEfcrDOZ
4NaQF/k3OjEM/om/1nW1yiUJ/kGrZrRw72LoBlVqxC/LSGASi1OJG/JiIc4ASE5b
zZGlv9FK85IImTU4ggaojxZDjZ5hSb1VxtZwbjv7GHtHDlmNG9myBjB1hjBMNalI
8ph7Z5INoeTKqcg5LcB0Zat9b4zYOcaMbNNl249MQrvGYYHamRp1185lAmGJQiCR
dVGskePR0ct3zv/uM0QHTAe/euYgFxpd9vy2OFiLzCiO+cEhC3i3lK8gRGlPSgRh
AtHbnvp1+FbEuSARdbHY8iTwKtUbVjAhzxYvVwwNtbgBP1NBelmSRYObXIjLOhgk
LnNcYYb32vCYSbB4zUmlO06IuQboCiduLQTZdxq12OU/z81me82nagbGNWrhcaQR
wkOfxcAjTthHA6YxKA+b2DLCTC+1neygmgXiURa+f8XB8lB3TOqm/YKlUC/ZUGgd
5F3oij8sTN/73ecnU5P8r36+dcqjqM+f6zl4JQu3UGURBAkgH9Mdc7D1biJUYgz6
UfL0fCUPa0kWzEisiL/QTTuvOmxN89Aehkv8EjE/RJ8iojTcxTm+0Y5QqIEmiWZB
fN/9EdBhukWRUETnqBZUzjgH0YxHOS56Y9AVA1DSVCukGWJRhcIomabTNkmGJb98
qw/D/rdyTih1k4FN6JlmL5FxWgZJWRTsIQCq7zO9l3KvlMW/dNI0k04fjuIHvEJY
y92PbENtw2d4CtHWo/19L3o14GiXEIj8fB1jOt32coCvqBcmmy3R5Gk5B+JJpMLl
V2VwW1LBKVxUJmAJZMseMipctrwa8tg4ESLb7AKo7iBk9022GEzyc+OBUoF8jbev
OW6LHLnOh0tHin4PTn6Bv33unTDvZASsE4iK5T6msy20nWd0Fb0qL5jm65B3f9Vf
snD4wigRmO8ci66WZ9Yh00pqOGSxcjZ4iZiRP1lgngBz9ZrxezOP94SUx0ZJTHH4
yFNNNqDq5WPv+hx1taycoyGHkYKPaePgcYph1S/ZED/XI82m2TGPB+ZtlXYJJWbe
U9AHNKciGqfUtTO6ErReuh/9dHqbXgzXOWzSgUxkLAACImvVTMXtcDIYbVf9mCxB
NwxCtEWvKymZl7eOK/jFcWrAMKN1hu/TKKA00jG/XepaXmajdschTrCa+v3/sXus
WXgQx6em/AE6njQpQ5i8hqV++8Mo9tojfrJ6i0oWz9XMHvRQZ7Ym2nGUtlWPvtbk
M8bY3KIWWO3Yp8Hy7xi5LzQypAda7rpsGjS09bR8yd1KztJboVnWPmxR5zjLQFu9
Ujn0y4BYF2selHHKsgGjL5vEcWCdxcGSABdTGiuNwlZev4WSNAFtfW3hV2i6p6Lg
miyFXDCPXtb2ALUOkZUfNAfwzeW5/cGaIu4H2ZrdD9vealA4inDbh9dPN65dXRRy
KCMMsykvTeCQGYtD14tzwfvZ+tVS2Wbs87QrrowwptSUj9gxc+0EKNDynqIx9Cvs
lqXtosZdjbVstni82xWuZV+g6pyzCyhCQKHOMbDeCFuRgkIAWqYSeiHlf4pdboEc
8TuXplCXjqtfJALYPZzRzQIlsJlLSaEftvqgoR+J+GivI6WJhW8Xld+zybEcjfX8
XgppCpAJhS0AIzbShHupIv/sLv+r+JGCVGf0pZRSFMHV7h61b5wkkBwrpyB5Z+E4
HsqwLtfxnk9ZFffJK9hcDSeW+ygUcaShxcZ8KfBQwq9uzvO7137V8q8s//iCc8eS
M+BA2VMpSBum2LHyExTqrTZjpID5T/hJeYQqVhCCbtpH1QwRnsbSnfSgviPvqO6o
TZxS6BOaRZxjJ7xRaq/fpBwxe5xQozyZYe5n4yPE8UZYTRaFCn5bcDpdnZGKJDeY
7NB0tb7IbbxCrfBSIR5Qu8GVaVUkkWZDl60zHlL6hUn2deqnzNgHfRDidyxGL02T
eXQlmUKX3yWQozogWW3aNdLqyURteo4St4k/mf46hYYVMAaoP0VFNfd6UYsSZpOL
dR+5CogQhieaJBgp7em/5VpfGEgUWJ/7nhQJP8iYHyKiJOx8b6MVO546KcrOs/NF
n3gviyfTtrnoCpriPtOp60uo/6SIHEYPTNrVaxjchS3CiiJVuaSS6o+ScR9INDfW
RRDmUEhSJxgY5u/JT9n4Oc5YSpkS4kGjxuD00Z/gXHA19hsReOVGwnKOgPvRrwMJ
5XSu+jkMBivlFybtYTTGPUrlSSBF3VFhStkYmxSPoIoxiJHAYnliIAM+y7bijWfC
pervtzIdUiqBtC6VdE+ITU5y+53R2vZZsmUPOUcpUfVtDK3q8gZjNUBN1tzvhK7R
9O0iGN2qozroQL7y6u+hqbmyFHkeP5kA2lavLFhWm41xhUbxaLL/O+Ff08BjE0Aj
+uYJ2z+XjslDDzMrQOuQL3OlbTuPu0rWuX9Gyop8e/AqxP4z5WascWDL8zkgyr52
FFlldwdwzTKoYm28KaIZB+uE6bjekjG8Es/pc094vjsG07+bBBhKrPML8moEbmBH
O+St7w1hG5KJ11K2Fs0qf2V+XNukT3jaZNJhdOLH8rC0GvGaSVjODLw1A10otIIK
iHvkSZb3Bz9Qwp1W3RCBVY9e9xEDUUGAFtCMYtR4+LN5rF7K4/Pekd7pVy8XkSZ4
IO0UE+dWkUnPJmUAK+o28jxSDa/QBaJxDAVhvRPm60mZtHSj8WFV0iPgH+Qo4wD2
BMPtbXf0FVAOzDNruWpexgGvr+KPZh4ntlc8C+G6IPNYiZo19zokJshlPRnOWNeV
6RoIA9THQ2IZsKGrWCRPuNRyID2GR89qlR9R41gSem6moV5qjb0BVbvlkQba9KsB
K40+5Q6KyaKYbiSyIYjSf5VNWlNcV/b7aJkKuNZiKbrnoO9jv/pouNGwJBdz2aDj
KvBl+qNZEdAa9xCIbXVUY2X6dqgkUdKT1SkrWmZqlssPVyT1wcuTKIjN4Q2uT2LK
y1I6hEgyVslOBQOzc+hyhCDU5KgR7XV1viTutFB7aSyPa6W3ngnVa3WHlKWRbhKt
tFeMwAnqyu4A6F/JA3lTEQU89aChVydCiK0k34C3Yv6hTbrF3tw6JRljSwHIyg3K
BtT6EpAb4XmQtOuHcIqdDpqDmz1MoE6e0c4QSFsV2mWL/tUJUpcpj1IFLNZYQ5Oy
iM/IoAV351GSioqOWAEWTktsLFBeMe87UR2IOTFT1tgxCiOXxzudOSv4XsQJ7R3O
2Dt4bwdAKPsmlKZD77CKXe+8/A1eheAkJQxZcRxQbyb/50r3zOp2Nqzz3HbRClrT
qA3XRk+RRkpDWMz8NHmHhwkrmUqSt/7F9GV2M1aRyhfy4dEKpAhggF2rbdZS91B1
k4xn2oSkyw14j6lHEO70Eyg7bznv7lkwylrwW2g0SnvLeATSTbsJ0Y3BlbYy6MMG
sIES7AZIATOL5Kpj9e0S1w6bRgrkNVsN/CO8hIiCXD4+AGulbcEiiyuKMqjMohhq
NJ9SqZQS7RkPJrYJKw2A4ZTlbNg/NTyx4SHWfM0MtQYiuCeEP+mOkWB2mE52rYg/
h+Tmhy41/Uv6PXBOLQGtfr7MLXqnBNi4i2jOvWjqEg4qIn+VBYBKiPHEKgrJl1vA
D9SUGGADh2Y9F2ENCCi6tIBGcRidcP+gI6NyoFn3rmPUtqqyD8259FpI4tpr+KFc
Twf7Gs4CbkCyw60N0vtwlee2EUjNax9xkajLB4n5Gh12MJSn3tIQWOez/GaIAuMX
bhMbDZIF6VNuQB9AypRCidj+f2WTd7GL/GCFurZdrdl//+1VKi4i6KkrAwxPOxWn
2szoOUFub2JeSYBRtN3X2x2OHydNK7KT0BaG8vRkcyP5aYBB5fZwq/ww0q93/Hg7
sKrxToSnhl3rvAXKNwke7tWebqHobqDv4GtIs6znns3+6jxbarL4tBgstLf1yys2
SsngWigUWFiBxuZu3wZqNK5M2insWPoYkhJzs8pCiI14POBfntzQIt7g7BCg/s1Q
bvglvSwHJoae4DQBYvH+b2xtITWXdy26O86/uFXNc3IrJgX/1aHdOYYe+akReTVM
CiStEQ/TZss3W+0G1cN1xi8Nn7EMNaKmqNEXFe0aLHVJOlRjCFPF+nIvoBA7A0GS
QR9sT3CYROorlU5umM9UH/Tr0VfGk6VutRfeMCIFeycjB6aHc7u4zVzLg6Y9fCgV
6AcThSWCx4UmIww3ZtShSFplZ47WpnoEXUVuf1lRZ9JvLzypG9VOystglR6KVHVp
KUuD3Vt7rP3OCl/XaEk9X3ULcD0I1aCW4cx6TZVTiZEe+0YMPwLjQ+1wyd8EslE0
gvWb/Q+QAKdWBfnLVmb2m9gnjCEHczUG9WKZLuBKUenTq/i61J4mIvagz7O685s4
CiSJsQm2zmVsCkbmzP50Euoh7i3RpJeSWC0uqk6M3B3t2oSNVHPWM7M/0x3jnmkk
0078eDzZopYKhlCLetCUXk3V+c1L7UB3/1VTXvQIcsdIAQbnwtUnvr0W7JJ+cYdF
MfcYsQ/WivR7TsdjIPPBvphtabK/UnWG6QSmgLy2ByoWSiiu+qoSuUSR/Dt1la3Q
4UYO5f15eXCW8kHvkqUhW8Ee/E8NFbX9w8UFpycZ+yMySac675/rj9XqOdzKAalC
65JpkeYUP3uRlIvpI0xQUlFvwoH7fRDqKNWQ92OUXQHMEKom1V8Ht8n/W7eM7zLn
CVFLngiinrWLvVVSjfcOGprx29f27H3/dh7UAMKzWZyL0HoJYe79pKvpsceAVCTT
mhIT3uyMpVX/Z43W9A4q0cYTvadGCpCCUpq1QKcJQK8SS3wXn+mwDypABn3FsWGf
`pragma protect end_protected
