// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:45 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pl//tqRDnuMVJOQjaO5dpM4+pP9IwVh5uKLkrscdUZEYXT16i5n0v/r6QAO+wQaf
Inm+fe5xV8b6XDP1dcp9MgMutOjCDGrxjMSUM/r2g5kcHzgNq6Z85Lshxnue1jyL
RVWTENYP6bcE/DDPb7Lp5BDK/ZAW1y+PCcXGgDcHfRw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15888)
GNzDo7+l8DHTGlLB/fvuA7mCKGtz1Tt3KxEzQqAi2S0wgk1UcCJ8XbnEXkWGrAbS
+7vroHZKHm/bFaz6TmGdJoGUrnb9dqO4EvLxfb4ubD7Aqo1hBumNEfUkY1zYDL03
2fn4yGLCWZSbP9p4vDjtfml739aor7iOepvoVxGofVxIjQQLYxEKPxgvvgdIQ4gs
F/F9vcnKqUEt6k5qS6iZJFTijsfEcHKL6trPFvbf/oeV+3mcgjGOo19d4Ovftfof
HygjkmuaeGL5EmlmMVnz4tY8mfXiXhTJ1h1Q/AYJDeHqAyJkCqMljTugXilENJBT
gkjXAM8bdzU+9cjNHEIeBNOjety0UkA/1gf+DeUgdkjoKJeWVEA6DlRjzJMqyEuG
seG0Mv7kTZuRVviRsvFoS4lJF8orXsCdcNSgV/dCgS98pDgJbjxuqQsUZKPGT4iu
PMb6zu1coKeMnfasDIRcE8/LRnPnmAotV7fzxEIo/CzzVNk76oURF6rKQiVzIqWf
SgUuhDTMbDDfqyw6inNM+FDWsVABX0aM0yQghwplUW6E2Iud4fg1ZETyG5Z89ohj
l05ikNfzSS+B8P0LO6lCaIrTloJYRpmTnGxFmg7B3xvKnsKuqtwPqQumhiaBMinX
QAb8LxLLhknpubwEYRx0D2xvGJVChVebF9Q0Ziyw0wzdcjjccgvXyb2ceSiincbw
ltptXmebSgfs4Cnp2JUR5ou80p+fITxG0kQflTICz/Siomv9Qh3d1/YfKpuTnvzT
hETyDhsM4zXBfWzYaV6P1RXFN0Bm5USmPCnk0sza7HT6IgWIzMmr9zASqwbPhrm0
3DQvzlN+wXcHML1kEAZOQmziToEEzL+8jcFdyzOLwfpnMbLxfchl3cC9c8IrpASO
gowguvz4yt6MDP1FSNqNMfAwUL09hZx+ayDgDnNE5gHnfTpgF8OFTzia6Pos40rM
tcZsaUaWtfXOdMUsmk9xrZS1zqU9gZwzNk8YnfQ+bqhnPkfM+SGf8CXeydevZItN
/4yg2ivLa6BgQUoDa/po2tO7mL8r+MsKqTC3BuC4ZsFLWHn/ZNVpVeh3K7wcWM0g
Bxx63Ryd5QDw5DeashaRnRRHbdvwXRP+zE8/GwRrDv9DWnrK6RtrAsJu4Wj2Y9jo
4IeAgJ1xIXiqmlTSFogu9+F5495l5nU66zerSBYAnNUTSmFo5vK8Ryn5/X9I2ztv
Ir/vCMwueI1OsAfV3Ocaz0bvZYyOmexl9s6r2jP/2atyy7yuWOKZgjoQz6E09fAF
XXHqT5HaUd0TlutXfEMTf6fCdS/JMjR+kVhz9aACDyXKaeAmqEdI/a4PFrfs8ape
aVTXN4Z4RwgzDa9NH4E7Jccq6SuBxL/cnhdq1ZgQx2IvqIROol6+HFdurGtRaNBA
zl6/P+KmatY2nmAtNCt/Zor85nRdPFvlci1cC2hIP3W/IjNQbJBYqwpuGXynKd6C
mVcWh/+yF+Q4eC4Tizvg0BNWFcSWL124q1WqzT2bSQFGsBdUIOUpLSxf1kZM4O0k
vfiFsCNnbB2D/04Fo7T+q63BFRqL2jbzkRTe46mFBauSFHM98AF36g9E16QkrVv8
t7Uvsjz7Bx7Fq0iPKGNo4k3K8vmlpoAykj1zhZxXpnVK9CkpubSh9/PWjiwOGAoR
JoVz1cKxuvoUPANWMBaCp+AzTRt3XzyJp0q4Q4BJAfYG/oBPxHtZ1OhGH7JBuA4+
yhZpBaiZ63PReQR2KcmwLiIACdwz9Tbqw6lkRpPYHGnvwjXCs70QdR+l5LE9ZIP8
KzG+gfK4fgJyvWcYqv2Ma7n0QhquVJjedVduPmmxHPIIh1rNnwaj6mKRLxFDxYLk
YM1bRkoLcVBCAgZFjWp5ZpEzJglFqcVUF+BIfaZV2IcWoO066Kx0Z0CHgpL2CMMl
WY/n8ol+KAxbwpTctDD0tOkGuqc2lCPjEs4xKYsqfMNXpIYCZZeXPka6gWdpJ5kE
kBPiAxhRIL62oLfvQCMUnO6PjgTQLY4xsukT+YBFdMGQpGNlmB5+bKLWH1LMda8k
bsIbfFRl3hc/Bm5UAKLpt2EJv0B9Mn/JYwJNkArUigl56kJ+t0B2xfNQV7nA1LpT
XD1+SOzXMdzKLx0IfSoq3S4NHQgALLKqyuIyOVvAn9pDgolPUZrxO0n+h2CUfkDl
hchr+a5JkrvDitLq+cqyPSVkxr76+uE9yFvSwDO/pmlCCsOeze/vQkZTgIYN4DTP
P957jYBonyP8mLzLe1I6KIv1U74f1GIuykJpJpuoMg/QPMIq+DOmnAOzDUoc716v
WhYj0BFveXpR085hddJkzv6TQVzOeEQgaj8LT1Gv8gVZ1VfVemao9ZPyvg0jcW7l
4bIq+CMXjUrspFxtCMt4Q1tjT8yps6feQlsxbGcjimYRpn7D0KvCVl+fAuJ8OeLI
PJJBytvJ9Z0349JOeWNLRkCj5BNcCUY1o1tOt6mK1gew43mfWfRruYAKSGehtz4q
8mD4YEHkGTVj7wTYSlwn+mqwa/3M84jewsWE4Jiuf4NjE2I3f5GAIh5o7QIQi9eH
KiMXcnw8K8qShqIm0YdZVhxyJVbX3M1tmZL7J99mjEPAvLQ6W12l3lnzGsk9uRXX
yvfQiUgkP3CuaJljwnvkCwQn7XZ++S64zUPAHwcOKYqQHhF4OM7lfj0AsRYG+4/x
Jztp2xvwxR73UUsxdgR7bacc5kR4mvb+lGr/qjgVota806nQyNTSmiK6giY4q5J1
WeFrtr//wR7kPCL68eOAhrx8g2IsK7Eii0FhkJEhxS7uxQAef3hm+cRRVGEmxeAW
ZTgXVJgS1OT1tLzlUSPylQ8ei7hVDkarvESfuA01+4R/k4Rn5sDr7mcQNXAsAqqU
rCFn/bpp5A11g4HBxx6IgLppKBTVNzz9o8QgCVY9yK8RqAXKyGoGRiEX+8GH40V7
vmPNq/gPO7xgGo+kco4AHY4xvYNGEfZtVMERrhhyOfSXNo4SrrMvdhb2erCs0iky
ho0quRi1vJ57Hf7fJR0MtjFXktf0+cL2ewjKaBIGBCXShjC6stSNaJm28wxBQwSU
U9Wbio+GEE7IXH6QFuzPkGJAv/8A4bl4zidVa23N2HsXLkoourdFNd68IopDLqTa
mugu5ZfPsyf58SU9Ma0+0XI/kdE7tmFXSpvJnrXJOtjm6smJl8ROVmyx3H++Pi9v
xfC9zbRSvJfM4YM48V76RVLpcJ+bAWv0E8haj52WGZZYAJyfbQDcrhdcW9exwd8x
xqOMjIdg/N6CFZkNy2zkxqN5PLJhyGCB57of76zAHtxCtR9sFXjReZ4qwq9sO4/N
EhJ/LkVYBNbJi/1+mG8i4tzZlU9s9ZpjRteNB9p1cIOMrPdetYeZYISglzPoShHq
KI0nZSuEXe2i0FLubkOuP7mTlA9KL6714Pi17TIzJzeTGRjir7v7ZwH1rl6gqlN4
YgzQMq9LWsWzq0SPxbBiKM6/6iDPyDCDOfyEXjieumLajOTfyDdqXb7Y7RoFoq2d
H94KTY9SxNGfBRmarbsXB+V8K5RaQNhx5YFksT69qGhSkKwmUW1YjQrsf0tPr9Wj
P6AZnDQ7zlGHQJfIh6Xz2v7DYox3eevpGTDwBVuFigXDCf530bfrCrulfg1IfejU
hThS0z87tFICIcWl/drW9SYU54Gn3G9lJcItoK8gETf6bdoMMwM3MbZJex+zie0/
/XUyofYMgefSyDQNnZmERYB43o8UjVESd9+s8ebTeYDGGNUtKMezzcFuWTONuSTG
/juWk1GtNmSWVhcuEtnKsaEVjG6aQAGTLcbskKqOr4ieXrP59a9abgmXl6VRIQUL
MNXMIUYXxxR5l7k5nq9G+sNWtAzq8RcghAkbmd5Xj76fJ7jFXCtnlU6+Wai+ve9U
jgG/c8NphYZ57Y1bIqM2Ph3CggI3aE+4XJh6ScY33+YfQjbPYQZ+rrvweEIF82Kq
y+CfQJKOhNr2WyrZGKjFN9VwNFzGYobxa7vRSY0IYE5OB5k9B+Bk1r0FMk/sxzjQ
/IhK4eBYwke9IfyWUfmfxQfeUsnqX47p2dOL/UvlfD41shrVg+uHE84fx+tLPt/7
hoi/dxDuwsM/eGTHu6sYywMap7OSK3Y+f/VAOs1gBCNOcSCed4Dc49ZmwBDi5cae
iOh7nHXhZIONgF6/ql2Dv1dq5GCACbdCGJma7fhSmVzF5Q396VdmSlnDFT/+mQJZ
0IjYwP/bbSjrw2cYrueLRdZ3JInqmEynaAmnd6yrdYr3rReG5LViqRE/12KwwGhI
b/8+HN4F/SDbyEEqhI4Ay725teog6wvNrb68U7Ei/MT6RGKgZXKzcmGXcB6gb4bu
SlLCjHJt3b+WyAM0zHkFOSiSdFG3PoLmngkpf6fT9lyeZyM5iB3OOMMOMNzRiSX0
H/le6emv7K+NWbK7KeVZbU0UQh/MGTwOkwacpFeU3gCW+MGkYuo6mzt90ha2fgAq
bPgouWQXRASjaDpKXS81mrrU5eKd7SwmAqIvzqweaqFvDq0ay40VUpB0FITg2tsv
fI4aH67orill83U3PATewF3Es1jCNx/CVa2iRC6L24ef5RAN1LqP4Ce19e4R+oG3
asxEvaZYe/FzAFByWbq1ahma0/KLxW8Phpwqb2zN4oWaq1tUzblOf3WUuSYUVTpU
0fhOxGgOrJ/eCWxW2Y497L48uAGkg9QPjwI1iNjfF+iR3QFMu4Al5Jal3L1y5nSr
/jvNQkWhcgx2Fko7OCDD58Y4Wc2C5kQj2aaL8D5QrLU+6D+uVFS4uEg4lv629fwD
o7ZpLimoVdzgYjtKy7fpQPAyBtCP3yZ2tB/n2cMbhKNetUusjxYWbn916Q1QhCfe
bhKB/mzh0qFXvgdHxHGSX7H4I2wkiJBzkSfJe3A8j5L3usomsYGhkFBQsGa8RrPJ
ZCdKiKopNhwkp8P8o8HyCS7mC/+TcGIj4kUf7OqM69VDB0V8BjmOQNPaanw8RhgD
XkDhVzbx216vGeu+VDCZNfM6+Im+rrLs/7I8eGLIGGcc+XR/KJkSiqjlVVZixFyK
ZD1z4A+znosWQfia0ylZmUXiN2SAdQpg1nDFtOyJrn1/BKpNhYRhR1vO6Te1dU4i
WZwkg7m1v0cIqUA5axUnt6Kp7KDPRuHBvEH0mpzTAhs3LKM/gs2+X6/UdNO5uKb2
Bdrw4TlTph11wHkNhycvnAvzx2kqtxkffM2FjngMGPsKMJkoKDsr1Smz+plU5jz0
4jMbj6l/FBeFoK1u/bUdq2uIW/XWRLHFp8pqswgPSPqoxZGzz2X9FHKNGw+60baa
fM8Gi/4l/PZQ2qbt1F0P/tYA1oW5JMWuCEO8usgI7FoiDyWpAu4+RmsKhBFzUGHj
Bu1O/3ezqpNdbrj4Dg2hfSbyIoMROeNKZUX6crHIOnuhSt5tvULSan5Up7wCAxPr
i54dMfwwufzs1+e+IuzhVLmhcYhA1JvTGUEGTXPHZAk1kKtK27INOokOuYUegdQJ
hFGtCmpmksQqaPzWbm2CKYesBrCyuaV2w8Pjs5BHNB8pGMMSdJv6SGKoiEj4asIF
pV9CVSL3duczyd834b39eFBofiaKL75e2x045uXxBnoNfKPG3jaJcASOvENu6iyx
tAXT6cLOdXugQFyl9fqZyKd1/c8IAk/IlcorHRQrsIN1cJmAZVR12P8W7geN6Mlm
PcKqX3SKhgcrQyMcXrc1qpgpMu1iZN4Cjaj2E6x0ERF+WNgnZw25aDZ7r8DOYbRT
nKWXmqiEVzIhh6WaXPOYsAay0FA5wBrXVF+JMvxpOq6ATL6K6i3wG31pT9nP5zBI
4yFjUGBQsaoU22nNr6hbtid7wM0xx/NhMosSV+sp0oD55oxWj8QzcjcSmTEx9jaz
B+F3lDTz2iFSCzSxcHSD4si4/+qtc4a/+MN7wHs8He67C1/r3VO5Z46nnJ+cmBaP
+lxq4JnRlx6eNTMPvL1bJ0iPJCnZxQwb8moly4E7EfWrgY2hLMFAN1j0W8x70J8P
weGo3yhLu7Eob8zP1gZMZmpH5nOvWukcrYd/RuV/b6jDhTAHRN+TMmDTUI5EsODc
t5hEzTNJ1i0vRCjpmH5IeY8njUp3sZtlssL/DelFuhTFekNHzV8Pp/l9BQODRpfV
1bw7+eYt11HFfQzCwgocxytVuqjK9a+E5MlkpiZ+p0X/vE6DAOEFaVRan2fkSp5+
FLbrhdFzY1vveM9Tv2/LPEVdIctHq5kPAfYOL3Cn92iM6RfNbwDyugjjzSFicUrC
QP1+rl1HnSURDwLB3H6dsL/A5TJKuoFI84M6uxYRSn4vznIDOLQ29sGjLgBgCE0a
KE4i3fR3/3DOK2SbuSbzWbDDLeeh+DH7S0msNC6sQOfbkYCeN9vRtDS+J7JiTZX2
RE6wX1ZJqpyAcrFMygraVXsAPIxsaEYn91rlY2GMJtqfC3R3p0jxgD2VKU86xmV2
Gb58+0rZaIIVbTP9tRQFO+iPdSIjUNzvw6Ea3GlWCGtbwxiOXTtWptzaaEI/QZhP
eebzBSevVRNnHrIqVRXvogzS5wkrT5wkyzBZSpeNnzGb3Aq0TaxqkO54b1IcDOME
owOiz+V3w/niuxVCfEOL9UHwd1uCNJw3D7v5gYD7X0SMxMk6sYGoYupqviM5SNpi
X3KrdcBfQtYsOCUdeXu7tPR0fR/K5EiUFGfthQ/fiPm9MnwebcrIH9+hxb7TojHB
ujQ6m9HSvyjgcqWi95gHk1Oa+z0EQWJ7ak9M9ctYXoseAn4LbZsJmaML4SIwD+34
pjixduRC/qy8l8YE+Srbm7Q1j66eXMljZMxG2+2MNa9TEDuiJcZZ5ViI6FH5WV6T
Yu/dUD5NxRZHVQZUxESal/WH4o1vLXRRheI75jhzi1JpAbHRFN4t8Z5dMD3Cp9w9
HyeDA/rS2l6OhxkJs8MmERT5CjjI7gW8ZKsmE8MU3OLTTwAckx0wVvRBApfGgzmx
s7u7pvONgiEZGk3cwYXhu3y720fwzLRwR0e1BqF9NuMo6lvujc8kzDcvyyWt2NNY
D9NdTuX+CoYbWvA+6n69VHXg7SvufI+1eK4EgmiVkm35QEaHIq+rXy3m+EV+9Tqf
aEc2UaEScC7S9FN6cQBM1GNLNtq9db2jgSOqqU1cnMhuG2biQtPkWVLFhDIGkXyJ
shdUB348UeEqaYM/sJ0GZvmvHseIceXwOg4qWFFBUcUCnR17/GBGLup9bkyfwbcC
hs//9seMEJhLAMhTzPKFvAzi3mg4ake8UWO1WNW+xAvNFnidekNFstluQNcOOJt+
XkNvC7YLRxqFCBhXoe10onXlRHF/QLDCJn0wqxZTPDsAHuf+Jnv3PskKeryRFb4z
AN+JIoM9rSxt2rkaZrRPenH2ZdicVwI9AxaT4vJ7fCiOwDQVPHQWtcpJyZeF47Fb
EFf3eLofaEYS3I7FY0Ig3ohSRGuWEd21SviTQf4C6IehZ97jtlh2VztOhBo7Sn3/
qKLTIRjGffp+x1cJRVi78DSO1Nmh+GCEsiAgZler87rn6DS1glh6SK1Pu1y69KKi
/D5cIk8o/nLB4Zl7e+5B3H0WwHXIIHPfxfVFE4/7Xx91xjFd8jrwuVn4ibRf6TV/
mMXh73TvyNnCynKjHbuIwlXR1q2skbENF45gcdrhcuWMg2xPH6Fe8oK1l6rKGfXa
4e8dI5kfpcvKpzic+wn+5Zf4XHkw6ulNOpE9olQjE+xI4wxHedDRONCAwbjYjZVI
mj6JzFcQ4owE8GW26Vx3TFNzGcugh8fmBOftaItyfZe96FfP3VLS0/FJMKUjRRlC
bl1OWzP6cRc6jc+9D1Ova6+2T3HD8XSUhs/7fCf+3VWmseE4qVjgt0XsXzV1G2eH
mK4K1hELSnOpyRSHPp8MzF35YhlSItAPwm2Yeep1OMnre+rbcfcxhkR+MNU7E9e0
yiMUPbAGxw3KIHtubtk9GlN4NlDDHgPzeONCgYC5wVA/HDnfOzOxFDNzQW9zoRQf
zSz3bZxCEhV4w+6rFfp6manhMe504eyDfhJGvaKzzdrnVpq1bYoyhd4Yz8V8N0/j
ycRbjm6A/pxtJVc5g/N6IGTVS19HGUfr6lIiUXqjKPDgeWheTvosS0PrEXQZMdiT
CHGYo0wirOEygAKp2HmCcnawT7CLqL7qhrlPBkKpcpl9pUDV7f+rgaiDet2pILIv
zeb1RIbY8ma9wVXtQ2K9dEoKV7N9U6DfqMWHD7GEeO2CAnuE9WGoFGDY+JzIwVNQ
3h3kK3pEb27M5nxCMcNhRGjgeAHFTZ3BMlJ8Ik28rYcav2HchC6LzGa1aJgmcOsx
Li79Hy0CcS3Xp+tFpi3GkKXXeIipOkIa5DO04F3rjfsHUvP+Nxu93EB91gAtL4lK
DNfKMWccqT4EABNyDFwSsbanbdgoFqunIDjxqKWlo7DgyVNdcl3ei4Ix7AIhy2fe
FfLSvRLTv4NRO9kFWcE5S9UDeX3fsmiTYU4cNd3VYGKxTdu5UjvqPPDoeaJESdG/
9CbMfgng+5o5wZp4DeYNHINm2FVEddXS5xx4avbUtna+uyFPdwAiYS5eLCW8swIA
H0nRF/lNbi6CiHQpsezosetDeAIQGqGA7oSQESKaBoDE3W2kPTF1d6Qdc0LK7xH9
pswyPzU4x68v504j/PngWnmpMqoM4vMbCsXE+/ro+oh+U5jZvhQApOR/H6G205Qp
6Nj4G5DG+HtruGi7M2nXKOz4BrAJbv+3aXcFuupcf+H2GF/tpga4I3wDZDNqd186
CPlqkkDE3lA6oYebOzGEb1Bt5eC3dJpC/i4jpXwZMCjF54iNzfJBXhrD+8dLt9GT
EYO1Wo4cFhBJi9+FRnaNUBV+QRxBpWOR+uZmzaGWdezvFJd5aWoctH0JrwqyL2TA
GHALrq2OmaBsHDt4ej1SwSiaSDsBqbz+O89Jb3qoPBIwomr//CFID/YDDBiTMjCw
eLQ7CZXvxMBQ/It8jjcOUqa9tNjroOpJvfUt8zIlFcrF0C71XsOO5GRuq8NMS2Av
yv/2lZ4wMe1RF9qmyKowNjb4EP5N1d2IHZVCI7bQyhKM9NdogrFewR8pJK5IYlVP
l8vtA1EeluZBXKY7naV2ga3N9UBUj0yFqKKXxxOs6U1h+dw2wlLQzFeY0qK9wRDh
rK0BkPx6wPbgHJZ0vpurLX4Omh/Y6jbfRc74VBEQJPNMhG+TVbH1xE7oXQFGnSTJ
1v51AVDcEsUQc3ZlIkh1lSmsjhNohENSlOf8isEqR5xT4rs1Xrw6+6BiYZyH7Wbj
lptz/RoLjZzI8yJJG3afwj9jf4izuuDJIVwi8Ue7SpsVV6V72IAulKIvGe+AAw/l
9TGz9ADYnhbmA1vPuRQTdQ/4QhYsoX15RLDG10whVEBvr9mtcrXc/fgK4AnQxzny
OsRlkSSRLXMN3gfrtkhuJv0NHd7YGZNoLAndLZkpRnBdDMDSd1y3iBa5n4wl7tBf
i9T48c/R3Z8xnxOE/HoFSEcB7RqLELVa6q1AX6tUMr/9Ke7RPOCp2fB2rdp+h8B6
IG35ndg/jKExXXPrEtZsQb2CN73E7I7rxBKeiZYtz4K5jwoMxHjojZJvuC+nPpW7
kL8LR1JbDVgOVe4teW+jKOkP+w2N8upwiLzDmiSerkaapN5+pq46U9yU6EMmkT8k
wcoIEsMjQQDEKwyGXxxPfK+21rd3aSIjLZFBngRmPDkAdRJtkDbTQAR5Uukz8sTR
SGBFTrdzlEGP5m4t53ft4chq7Lo1XdVHTzMUGQsZlI56oKXX0X6Fs2iwwK3y8XER
3iD7ST895Y10jPb+Cdj0f+yhGoliWTrJSEpEMCmh2XmW3xKGhzK8HwE7zxZvxMqM
rgAb0R1/leoLm7jrnDajRv/3iAgIbUMKqMYaEn/N92MbWvHAhcE7zNktBx0Lluzl
j9WyuWu382dJxXFU4kXBjRwjI0hR3DfJ2mVqJAw0queTjAov80NEtOmFGkG9l5Bn
o1b/OqQbxjEMkUUTg44EwHwokyWxB58vN7icUt6wrZmXTW4E4Y8Z+nTP29iDOJJg
eoI8LFg17sn0rtph4iqp/cdONazZ9/IC5sukeuotVdNIa2b1aDLXy6eJBkaOB3oj
JMMhGUOPwV5/anXiCnWjixLYwW7OZ0hy1EYEiLMAUAxoQ7kC9mLLEN7U6uIFLjFW
S0t80ZjGBGpn6WcmqmuUIYY0bcpwtSB2ZTqWp1jwtWU0LAzjOQcbqtRkP5IujIul
U9aHfxbC6nu3sf7yeAthri8evHKIHePy/byFFkIGBzrX5lc/3QxNJd2rsc6yEOi+
GBUuyx6YY3eEItmeUj3Gg8qYORa2wlVAi6qGcR+8Jk7tlJ9enyWZIE/ycTQcg0QL
SeYQt0bw5wfE+f/eqRXPfbfG0ZRhJBL+4gODv8kYgOf+xcz2cgCxz4X8YQvvs/oa
bsuoQAoT+s7AuDTY5F0EEjo2O8NtTP+9KETrT/r09+V2805PFS94midWHraG3ood
OYe9rI3zBuchrcAW8uNDLhRqSkVOjG3/TAX09i/z47xhK7mA/zN7PmHXRzvRzN0Y
y0LwAoLD3GARvsWXCN+N4NmETp53UkWezmH8KMrak+G10T7Kqa6k2mV09lHjzAuZ
3R5XXxSXyQ24yn+KgziVsef5fXN5UmCmAsSJ6fZPhd2FHAQKHvfltIT8d4RCzyW5
wE20M2XAGYZzdyL+MYwIBvGJipRMtexDunGiAvg/soC5P2+6AMrQtFyYRZzxCJPb
wZkTQ1Fv03tVB0TI8DUUHKqX7LxR4Xj9q2Rp4aLDK2n9vOTZxhlaP35c5ymTFnw+
pGNX4G/HhmzOtvipRZe6ggRN1iUJstisUk5c1hULcZAO6uxVLv33VwVjub84wqqW
wvIWiVXt6/rN6128UxaqC2hi7G40o7ti2hKm80z8uLcwac94fViZ+g/9e5R4pE7t
1b7JCrNgII1i4yB+qHYNdJM9h6ypUyXIQoU+cgsAT74AnWHDDQ0ToUqICmoje8q4
xC+Tpu9RXYutKARIJCvvuZK6RCUQRuKsBYOkU95UaPV/nHQpCZ714Qrh9uaD923Q
yRgaouRXS/e6BiDwiSJs5kVMQxd5ZCnP064lrQIq7uBrFyAMeCEvVq0vdfWog9Lk
VoutGsHMmg+2FmcNx8RCwtE9yixcOyJUEkuAf0pV0Z8qBYfBtPAg4NW4Sd2hy4L3
W7KC+ciU3iLYbEoPkFvSyA0LImVg8Ou5GdOd39peTD9OvgFG5nSpbOAQCW8cPzbH
FoBnlwff6VG+ecISFyJqyZgPuTkHtZeiPJj/OLFI5AIjRPEmpMVDBRUlRyzL68sr
pPO5dFD82R6xyR3HQjgXKbd4Roil31B+IS58V6l2Vs99Ke2K+6oX/pYa4KbAns2S
6LVkn+ENJb8Rc9yEBPs+8NCv0pjJZP5mTW5JlJ/DUU8dLot66oQgzuTa/4SWT1jP
yrVRL1pjNjvBdOuXh9sX3HyKTnK9uJ+c801U0GY/E0h9vf+U719OZmFzwNeikmV6
DrT9Fp3Vi9sMSO0AeocidN0VzNlUROXt4B31eFUiDKrHmygHUGgao+SL4HDDZJ10
Y3sCMNUTuqLfiz7sU1zwOJTe/45da/EA1LsuIJK5uySDS2O4JuISOt/mHYBkwIKp
lVcku+Ys8WL+jMjUr5N6/cNG40R0kEsXD90nYjX4v/PyISrMEdU5xfzFthTPLf0S
71YLclMP7eOXAqTO1rf/jLZcWYyIRJ85pik4eo67CmhaTkAjBlNg6XWCaJzetMwQ
n3uWH2U9nKeBASI63/SF3ugsiEuykyZrzMx3HPRU4D2jJkuc7vOfpt0C7v/Z9ZnR
aOTw5h/kpUoaOB3FTk1N3sAISQUobRIs1uR0GRJmzLfoC8kR8XCn6YC6Pkdk5ewF
4D5Si+eous2HgWoKTsxYe0tdeS1BhF50HI5GD4VRO0Dyix9DJFrSuofszjp51q0Z
VZpqx+1vNyrjazsnl+Sbzza4W35k9uLVvlabKZ3eQCHeZDZ/fkE/NIBw6rOXV7ii
xU9XmZcfWhosdmOCPURteW9T95Pzy8BLz1QcQmdthBbwN2cAjlE7b/Tiwe9gQFZd
FRnJ/izbA3UhEnRU9Yvg3ESKJ8kYFB9d4TlAgTehub8OsmNq/Co3Fnnbfm+lh5Gy
AB3r1WF7cbvjOkvp554D8p9hSCXYnc3Xxg3OIY1zNCXvwJJQ+ahLkLBqgjrslIA9
+tJ8AvnxM21OukW6GTer6NnxUH5kAWv9lemgdYbhRGgUR+ImHu4PKAEEYPLf8tr5
AJ+iimvPyOKFkrXGlYFXdNkJU6awguJ/Hw1uYy6UkO0AJrZV92HeVwPmMt0/xg+s
cfpQouBiUp+k1lma+jw4lUjW3nVWLS7rNVlmzwiRkf0zmblv3ByX1fapYS4nO5Fs
XX+bFn9KUyNZDhAUI+ejOrdiAByl1cciQGLEgRJ+VzDCAAklkzXjPkpJuMF9ebHc
BeoQ5TvSWGFr98tCpbS7RqzqYquBP2UkIPqLZbl5fb0lqzYDzb2h05XVu+eaH2lJ
6fHPD7Vvj2QBt/g+sZhbylt9Ysc/moEJ0TEhl1pH6qOPGNN2IrYxAE0h9P2/T9qF
JRM7tRWvXtdjRwaptsagiqaz4O5EXpRWSam60jcHc/0UT2FeEFgpNG8nBCjgkyxb
RwqQgeRGuho3XAtHftBBSkhWAa+Mlb9FqPeVjIMXa3zQGLGivY7PccskDPg4xAV4
6lMYs3/b7bTotbsKuGQCk9ovRAHcecCOHZ/vWC7yDA9RMJ9z8hsS1OscNDY+joc+
2MqX/rIMB78BKLvCD97OUUwkfNGpVRu/bNX2ysMq50DHnOfO1aWiZMoUxIUClBF1
inJIMVidMCWkspF/c4Joq8YiA6/LeY9DFDRHlFl6jaQjDsnpwNo6JgtUiUfL6wXN
S4doHt6NrIMT4qnZILIFH9TfPCnsX1OPp02DJ30qr8E5JXn4kJhYEQHJrDAkXaOg
hP7/wAhRZujJ/VEZzrLsCa4o7s0667W9Q3Z7wRif+61YDOAgM9jpq4Pcm+Ujtpo4
2caXbdtSbf4ryjPmBnB7bAuR/q9CLKs8hUcBLnv1gAtBnPAa6Bv/kKMbE/Iu+f2h
eVI1mgbDwcYI8afZJyEXHv9mZzXfOdvHnATJAQMsX8p5ccP51QIVyGxdY+dCC8Cl
DtZXz1GVv5LOJB5tknv03dmaa/MemBXqXFUX/QN11worU8q0qFvCKpgHjaUtmxU7
qIgkQ08bblTL8Wnw+O4MvCGgFOALNU2dQQKY1jS0+IWy8ZCdEJLtHJFTvV7WQtlm
vLK2cySDFoTDqmF/UF6ZLTfwvLrBfaP05FYspVZOas3lHbNVc64Gwmfz0HzPbnKv
7QI88EFJ9QYHzFdYLFXxlpw9JG+WMP9u2XOd4c0vsWhn/iA+WcY6D6vCpSc+c3z/
PpE9tepB90CeYcSdklanVXNfEKlc0CgbhXjgqgBKZeQwLHFDZ4NP6E43F2745JZ/
xkE10D25IuRUF2h9xLX5Py+JhKC7kfUZEdQJ6DbYjMWrQd7LVE/BCyex/MsfLcM/
5oZlkItSbJ4PB9uV2jKWZqfmF8HIGV/EJ2GvT7Jd7T2oMOrg6+S51hKhxTHx5smV
bujVHz/VQH/8PE9DxokLqBEmTtymXeKKIp78Dj7InRJ2QaQF+uvR1kZxizzv3YhV
MVMkXpVxrBhQxcWYMSJaO3Z5mrtSG1djeOARwoXNFpkyn4cgzgywknhGxzfmTDB0
fkNzW1eRTlJjd/WPkzlyt3NN+5NllpF0JO/wFSaxS6bRvIFjU87xDnUerAzOG2nT
V2lmK911wNobLV4eRNysO2m0WJputVEoVdNSq8XthrUV5fjHrCV17ci/PvfM7kii
OoPCGwN7et6/wM0cfAN5UaiDSqzjKLpPcZYTCesMm+7CGHjG87yg4pjaC7mH9PfC
aCVSYONxYhSLvXrCxqpt8281L87j8ECMx0Ju/u8RxUx1n/IF07yjucEMsSKTLb9V
lakmYLZ0z++IzLb3Y+8VzhFqow/euIc7D5jWjV6uv6lrH8x+lOMqVcE2YuDuNSIs
gy5Y0tXLmdhXswq4VIrxQPLGIlQb/j1YxE//dnvL41SjDFgbUIItwCJw7r8HlqRX
2CESVTdGESbj9woFwhlmw5Ym/RmRlaMODPbCAhFtz+qO4jff+aonTCkdTge1GDXp
CPGeTFZq5CNkioYT2bjduFGUssV1YenegC5ywVQ60gSFRTehGHEpHYF3WXcHMqcS
lWXoM17pFqFbG+5H15wjFuKxrNIo3RbMbSxde42ADFmvhfLDTtSwEhoKAYesqIpB
HFluwOCe0v0Egt2jgrWYtZKUi2nR3ye30LowdvK4mwUPq6PNPQbwBsBP7L+e6bJn
YNL04U+K9mlrKY/hlSbWHYg9dT0TaoMO3Crxr8Qch4975TEMI+0eU1x2zAQ9lE9A
Ym0FfK6AORydmOC5ztBp48RxHprttuH3Tz79VFO8vJbat/jq/pdrEzw/1pY5FnoY
L2YAL/mlF1kyozTN08xEIaWkC5fqYMaeXnBdwhzxBgGCssvmvt7wBNi1usFqLWik
rooUc/bHvpCFCM79GChbRf8bP8t3eGMTjXJD1wyD4sMWuBvof+qD12BMu7SvWs/l
aeBQ55c8LpakzMbf8iVJ23NxrQko6jPgFEoQggFyj+mZyL1ejCnEC4nCB8XRcoem
Wbf1mro4HTb/r5gpaTvXW+jGxhVvYhOXKBdW77OtjHwZPnJTxbgehKtcmSS9MO0h
AVEFXRwUailhgPJfteoqnQF/EYykgsDFnK9uarBFjLIL2cICkkDRRDjD38i27TIl
Y3kv7fhmao9Vry0awv6CY000yaAzI2hPVQ8ucBYGsuGI2BWbqiFtHCjei5UnPGHW
a+qswlxKMqZGCjKaPU1PFp7KLOMN+UYqTjJTuR8BZi8YHEKS26OE3YP5H2VBYLbt
tmEwaVttWtv13jfFvgUYnUCc0Whdhvax7GbdqLQSUrOxfOwecepxQTDHy6CbFrjM
2Cujy75UDNGHEw5SndvZrtGFqMATc65oENYi9RwW9KVRrvQWYoKjGHCiGwMapjq/
IoamVqX7nAcP1vuLBU1aNNa47YnNRvYeV6AqLz5aELY46ngKDZlMqXZj4l82K1OO
mfsdM4DJla+Oy0nWQ091NxdAZ3V8mNW81UKPDCEig1Uk8l4Cvy5A4bgTwRkcJc59
RQm8XoLra1tpCgZuGzm02jaA5cZZmYbIekUouxYxwbofj/oqMIbfM9KDS9TsPMFX
/RrgZbzs3YBsdUS3vu/UchJxuRSYqfX/AMgaH/NlpH3MZ2Mi+h7hO/uDk+HS6S1K
LnIknpwf2wSDh2whff3STYxL8KJYCTp7+sRpA25Nl1TPWSd19K/yooYyD9mtGXcP
qIa7yS0h2N9ODskqKIInKRa+vE+tY68onzhMvdZfRieQ2pgvoeOHZj2hlejHCx86
VBcw/FZAeB7EFkAv2WL1PRcctbx6K6oO3DJj1+Brsua3rFvNutluca7Hksa/OiZX
Wfflp016xhJ0ve3GOjCNBELrk7n5aSCYrATFmpVbe3f2Dxllqcz1l0ke92D1nnTp
UBtf8qPp7hyRnxxjaddJNw1SAJdkibnRSfZ3IYtrIcdOveK8REsKsuMqbPYUzmhY
tAJDJd0Phc2McwCeBqluJkyOir1c9VXllRlmGRIPfnWQqdVMNK//LfMcLYfw4/e0
f3/vuQ61tgWb3EaKr+SzFZe94JcVEzoa0GzlM0xR1woWLYHdC182C+9vtOLyiJx0
XJxYhmcnza81Z/yusYPE/6gt7Lx/2cN4V9mcbgyE4XKE4s5z8F5vbfifiHr24Qxu
eN/gNdhSkgUo7awpzPBwwfDwwqXR4vuwFjtJOXRFZQdo+8tCfZdD9BCAiGHKwXWX
3I9Eex6Yyh3yADR6nXPAqO2ph5OnO1+hqyFB6OrTNLpFwpA8MXtGecLzsKJCtu3u
b1TYZmHq5GotOimQM6r8CoVxt3g9apj9qwLPTOagHscyotzkzzk9dHptT9uLcWvg
K95nFyIrqu88RCvMqjuJ8xTtAFumUSRlzJCNfilp9RaxeqCvd1YnSL6eFwPQ7Cga
cHHKuwJjuKP8VmrUaTPib+93p3SrfHTZV8t7bL0K522MprjuluPO2jVYmon+8hKh
e1KB/Q2XVL/EXAKylTVbV/x09NPqrttB84e0df47jg8FePgKsxX/lVhXhLG0QU6K
BK4e6ek6zYLTJGuk2u6E3VcdrTMtofnMQVVVBiNNFoOePpD7M+5JiiF08+kYITK0
Xguq1qOKLo9SM4gixKKuiAK0DWXSDvb59AZfY84Rbkm/0v+V48FI5wUdVeiFYnix
6JxQiVx6ShVLGUklBFlWhCEvmpVn4N0sUDDZKQA/Arz/7sTucd5Bj1a00GrtsN2i
87GxKpyCYxL1+e5UmjfgmispBLIjXIrssURMzrEIiFTCquvJ7nL/kYL/funsaWxl
LsB/i+4vpZnWGPD60HZSe27Csiz+RPK0w4b7uJmcNUgVu2SgLKjRs5xz2XpdGBvV
GMNk/ArRHrAUQR85w9IzZZ3oqFLBblnglvx9Qj+pLyCZvgQGbCrAP5npJif5wbHO
R5S41FabkDJiMpfVGmuLrJqH1mdlVfL0abucpLxKo6qN49pm4wR0LwrxO7j8UUJI
UCG5x5JQk+pgClpcBjuBzMcLwkW2KHuiHM6F7tRkDtSrxaMctaAOmYXEXCyIUYYi
FdBH0xbZh0WRyj6niZ56/4aSODDh/byClwtZiPqiEXnTGxYDP+3oIOhWu82iSMXo
xuUkpT14y8Y52KPlmZOdfZ4s4BU5WWxxjPb5z54j18Hr28FSW630Hnbj8h64cc7C
KuqXen5Jr4POeRAJUFhpIyy9gi3/BTENPOnztu/UcYKFdCcmzh25LAqOB6TfWnCx
OPFjSDMCCybk53+F02HaW19dI3tlMXmpwMJm2P2ftCThFg2hEqeVuHKSqf/hNwki
IbNdZscEHY2oJXgxHe5gAlQ2tBPUOxpDa5lKnrbQbDA8SZXIT0xNkvfaVrNNE1fh
VEyAFHpDVi2MWwwdBsrY/Hn0ecgFypOoCQ4ZAnRUS/MX8SfG8hErdPkH0pjYZ6gW
Huq8YV48gBHlg1NZ6xTHEtlCIcEXsOimM2ziVHCJ85Y+tWq7FgXzj3o/MkS5rVS9
a2HBxJCxActjiV4018yDysGrpRY/jUmA3AfIsOF0MJRSL7PuBU/vXxAb6OFTRB0b
QC2nP8mIqDk9jOUztreIvuHA+UimhWIMjgaOkElI9hdx4TSrRjQ0M+sni3RKviPE
VuGd4RahvTcACSzcYNAugI0vm2ndpGba4+GtCl2cZH8BLeQw7Lp+NTKLzE8wqCr/
e1l3j6hRZScIK1uYhwEOvGlOQFwsSluFTYouLK/E1zpGSfk7l+5Dxwu9rC2AYC2c
zd8dwEeDbU9Dfy5/Pk/Fv6uurJf+zSZe5o+CUZM3VUWSBesGsJstnNReTsGPgz9s
ffrq/Xv8VqCWTgiOQaILrfRx+jTrYVl7w+fuow4tvkN4yS7pUsOtxPQ2xWO0Wxi3
ebOlKIjYhFyWdJivYIu6e3+/PUhR0A60yHR+YsK/ebmpCwo1zUhwL97SJNTdFXA1
SLN+kW2BAnPmFikberrF+rnqE1cbkiefsBI4pJ3T9aXrx4PVqCbVGoGGlMmOku1T
w5YaZAjnip3Z/VZmZc0urTXUBMLfps0h4U+1rL9JzcS7wv4/fzUzsjTqsojvQTto
3qLgsSyvGVMNYbVncU0qKtBvIBWY8gXIJNM1f3pqsaUqNtkNVwiqfmfphw25GOp9
lPud+/Pj2fk3jg4CjLZ7LcA/TPvgzkHFoZ560ud8ii5YYy4GE9PnbMWu/+19R3kf
Y69cL6xnKJDZwy8rm0/kWjeKuXZgPvRvHiHluSawEXcNPF3r29p1dEEW8Tz6wUmb
8h7fd4b8U6Dsnff4abvBqY4LMuGDqwEbV6wpzpNdqscvCZ84LeNcrdEBB8E1pJNy
KpHNpIEmuuR+FcnWg58cgcmOVLQoDzy6IzjLkwnO5h19khNBRj+u61/3keiU9Ff+
AP7c7hg/mAna+eBHGtxFV4h8p2r8ae4UYIbMKPZUyOE02g9Cyo8tFt/R+fH/PNHd
EZUH3NhyBYXSsDjM/cObUFACIgX36sMBeFPVn9aVNyUoBjmwu69ej/0bFrMoly0B
ab/8oc1ryGpFWIx+wWNyspno1zexsrIVbrFg0Gyi+5Ht6/TMiH4BbcLDWthq3ZkY
IlyrER59L5WIwcIn8c4hyEn7otbXFDlYiU7sruzUI+vs4DP3iWi5bY9NVZ0q5+zu
6BcxTHCxzJRILKsAuk/UrdGDitHn33x16Rxey0CNQQWpa/zwEmDgkkb2F4HewIm8
Y2E1+OKj8vSwopvEU5TlhnD1LsBJop4SfeuHuAalbbCl4wyD2RXBtTVngmzwdYkK
8lA3HiciFdYrFS8Jq2ItvfrJgrJ7oJDvB/X9S71St8hAO35z8Zc5OED7DEMAlvsx
QuTnzGY9KKKdQhalxXe69TG2//adbn2XtGNkFOkIW0CkdTf+BcX3owL0W7qHNiQQ
EtxiXwPjUVqbFcRUwUbKWtUXTwGhssjlSuGc9/bC0UFeDF5epc8oo/Svk/Ot3y31
mjc4r4O7PYVVe7hDtAEHvCJWsoUsIr8R4LoaUYPJtNbv3Np97wWJ2O4OAMc4O3e1
AeEouWlwTIw8IWdBCx9xnrDAsYIRNnT9mUBaxe7sfKky0JMoOOuSLGVsp86506w5
uXkKFozZHWqUwkj2LiYV135qGNFHW2+zd42NUL68G6iRCMJmiYTg6D/m6XXUOp/H
M/qJls+gbQcy+lpeq0jRR/eOT/Dp/YrnA/DkF0maBEaY3RUqUKO1cByLeT4CLRqw
HDhu75JUS/2SLBnUdSTMzXl3qXdGbYnt2+B4HBM2g+txYkESdTT0B+wxN81kLK6h
FR8ew79Yd/EqVv5BJ8zHWbd+6DpyFuFNV6dpburxN9wg0tCoMhx+qnQmk32uVJzW
P010CNrPj3WEBwzed7YdPARjsaOKZGyzfuJsqMrvpMQuUzrBoDkVUOblJR+7UT1p
bLCRP1xxKyazVlmkKtV7DTo1CkE8K/eJzPaQRhkCiAcDMsYvLjgkI6D1N219oTnG
B9pAJ0Ui590yZwf/PaeNfW9zWz/SD0pW9L0Z06KSHVp9f7MKm69Bmu26XhGGnrCg
Vi2UGD4U1RabOegrgaJbTCB9fuFFYGsk8kLCzo5opTYzHCv0l5urlle1pjb463Uz
EYh5vhxdZf0dIP+nD5Qsde9IXRcHXh9WP9B/xWLF+R+SPrePaU7sHWfu73UL/beA
V03qHHqeHRhIRmnM0up3t9XJ6Oc0vP9emgTXbaBr/VIneOZSE564UDiR3n4BOuNJ
T2P6vRY3hJ68fYuAsrDb6y1UYDAOh4FMyflB61s3dqylFT7dqOnoyrlK5E+9yh/m
pUDysYNmv0a1+QiaQksIFL88ZpUTDlq2xRzSZdBI6cUyJLWRxGpLaj7GqRpqPXuJ
aaP8s6v4fyosIfL40D3qyYKXNRnN//zVOtSIQnUIJX/kh02w7NXnefj/raIlwNLU
dYjYbH3dHsQBhyiwose8v6j+htNVI7K8EbPWfbd40v0CGZ+qeJqQL491cqx84SlF
95lwYFCtGOeJ5Bf9AZZR1Gdg2MbAri59GsLlHbq5N1gu2HqiKzqscdn9G8D4H3GV
6XkGH4le34URASFZSNqjeI+OE5sutEDh+nUStLRTSQ4FlRztv+q1w4HE7pwkD6Qu
einFJKd6mpX/SuKYWK7mBzy6AXaFScH3U/nvM4Vm1IHm2KlKVh/4IAlGL2wKbdSD
Y97jDssYquh2fnhcQhRoYofCkpU2q96Na+XAlECyNGauiB0X4Ry9CJ2WtUiDNd2u
PlqEPVaxVyl9liHbKEIoh1nDTOnwdP92RuRfzYXsPOrfBJGaNvgXvbmPHqI/6Iv7
Hd/f8vAiJ7VVHwYX8DSjJhkMCHK4SIWWK8PGbsH50hV3MkVnYx3sNdP8XOahUFNd
60Z3O4vbQpLxF5y7NBJFJ0bCf/eP6DvzZ/KJ1whnXpa/5Pese8H2ilIrbuBoofLc
iIMg/Q0txwU/0jcXaMvrffxgn1uQjeexcKa8AxTMxL+vBpoHRyTMdH8vPjoIUEtS
oPJatXZbiAuAZ5wJJYwyootpT+sGWhnHIjFe8+WO0B1TjIzgf17BRyydEkKHkkdd
zAHOG0Tb7sNjGrnJkAAEWjyavMePdGu+ftDVWdK2YxsDXqMIfQWZDnGtctQiA3rl
hBytbqWuzSDiA6oRAjZkzq51vd88VXdyxt485q8bvjq+fdC5O6ZU7fxBLMCF/eCV
r5Ux5vTTCyxvwax8Qn3w8K+8kH7CHiM0WSuwxaT3wApMHDLhZNExu15pyzCIbynm
pEQNZC9EZkj8GHU+Jm/dpmQYaRB5HIHcSq/YfizjGT0Y5GmyKe19O32tu4YmNMzC
qvj8xp0/O7P36ndJ22X3ZuxS5wMwzXv77Z5YLMNGWxBnSpo1fWb1df86bQm3M8nb
L0Ei5YN3blUm5OOP9vzPs44viwnrt4LsiII2dsinF0hWOczFfsDuWccD3qJ6p3w+
25XS5z83yJrO7QWY5hg9ZW6amA/Ux/KWrvcQ4hl6ZjW9DsfaPsrNLU0eA63gur4X
1sOrPn6w9GO0AVZF6psj6goWuTms/31TYLVyKV+qXB3v0dZrU2Z+i+Hm1qVL9pFM
TkmGiHjYAUOHYQ3O/aU1aCXdE3I9dGYYki5VzDrfB0YAFzSQ5K987eoIcfANxw27
jPxZyDq936iRzf4O6tjbXdeEfgD+PEczLbdRgJ14eGBrfEHlzuiQ+8Z9zfPAI1K3
9fQZThbIWQTPMYWWu80DV75Lwn0wFV8iJxqK7v9JKsRaKcXQCoZ6yqbIlfBKO+pK
xu8MQvFNvNC/q78YNI2ytQYqU8mv1DSY/yDyJROonS65bUedtED6cwKxIrh/YRYj
IY++JYlHM/wohf8ZvfJIxOxLKJrRnJQuQcgFWtiOQlVupDBcW3FGOjuw8xqS2xMn
+JAMmDtY44+yGh6R+0W4ozWrs+EjVuhosRotN/Nk/oPpT1v4UzKei61s5bCu2nW5
`pragma protect end_protected
