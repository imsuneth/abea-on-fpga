// pcie_de_gen1_x8_ast128_tb.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module pcie_de_gen1_x8_ast128_tb (
	);

	wire         pcie_de_gen1_x8_ast128_inst_clk_bfm_clk_clk;         // pcie_de_gen1_x8_ast128_inst_clk_bfm:clk -> [pcie_de_gen1_x8_ast128_inst:clk_clk, pcie_de_gen1_x8_ast128_inst_reset_bfm:clk]
	wire         dut_pcie_tb_refclk_clk;                              // DUT_pcie_tb:refclk -> pcie_de_gen1_x8_ast128_inst:refclk_clk
	wire  [31:0] dut_pcie_tb_hip_ctrl_test_in;                        // DUT_pcie_tb:test_in -> pcie_de_gen1_x8_ast128_inst:hip_ctrl_test_in
	wire         dut_pcie_tb_hip_ctrl_simu_mode_pipe;                 // DUT_pcie_tb:simu_mode_pipe -> pcie_de_gen1_x8_ast128_inst:hip_ctrl_simu_mode_pipe
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata5;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata5 -> DUT_pcie_tb:txdata5
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata4;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata4 -> DUT_pcie_tb:txdata4
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata3;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata3 -> DUT_pcie_tb:txdata3
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata2;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata2 -> DUT_pcie_tb:txdata2
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata1;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata1 -> DUT_pcie_tb:txdata1
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata0;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata0 -> DUT_pcie_tb:txdata0
	wire         dut_pcie_tb_hip_pipe_rxelecidle7;                    // DUT_pcie_tb:rxelecidle7 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity4;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity4 -> DUT_pcie_tb:rxpolarity4
	wire         dut_pcie_tb_hip_pipe_rxelecidle6;                    // DUT_pcie_tb:rxelecidle6 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity5;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity5 -> DUT_pcie_tb:rxpolarity5
	wire         dut_pcie_tb_hip_pipe_rxelecidle5;                    // DUT_pcie_tb:rxelecidle5 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity2;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity2 -> DUT_pcie_tb:rxpolarity2
	wire         dut_pcie_tb_hip_pipe_rxelecidle4;                    // DUT_pcie_tb:rxelecidle4 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle4
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity3;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity3 -> DUT_pcie_tb:rxpolarity3
	wire         dut_pcie_tb_hip_pipe_rxelecidle3;                    // DUT_pcie_tb:rxelecidle3 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle3
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity0;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity0 -> DUT_pcie_tb:rxpolarity0
	wire         dut_pcie_tb_hip_pipe_rxelecidle2;                    // DUT_pcie_tb:rxelecidle2 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle2
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity1;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity1 -> DUT_pcie_tb:rxpolarity1
	wire         dut_pcie_tb_hip_pipe_rxelecidle1;                    // DUT_pcie_tb:rxelecidle1 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle1
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata7;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata7 -> DUT_pcie_tb:txdata7
	wire         dut_pcie_tb_hip_pipe_rxelecidle0;                    // DUT_pcie_tb:rxelecidle0 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxelecidle0
	wire   [7:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata6;        // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdata6 -> DUT_pcie_tb:txdata6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl0;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl0 -> DUT_pcie_tb:txcompl0
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl4;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl4 -> DUT_pcie_tb:txcompl4
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph7;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph7 -> DUT_pcie_tb:txdeemph7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl3;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl3 -> DUT_pcie_tb:txcompl3
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl2;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl2 -> DUT_pcie_tb:txcompl2
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph5;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph5 -> DUT_pcie_tb:txdeemph5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl1;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl1 -> DUT_pcie_tb:txcompl1
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph6;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph6 -> DUT_pcie_tb:txdeemph6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl7;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl7 -> DUT_pcie_tb:txcompl7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl6;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl6 -> DUT_pcie_tb:txcompl6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl5;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txcompl5 -> DUT_pcie_tb:txcompl5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph0;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph0 -> DUT_pcie_tb:txdeemph0
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph3;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph3 -> DUT_pcie_tb:txdeemph3
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph4;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph4 -> DUT_pcie_tb:txdeemph4
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph1;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph1 -> DUT_pcie_tb:txdeemph1
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph2;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdeemph2 -> DUT_pcie_tb:txdeemph2
	wire         dut_pcie_tb_hip_pipe_sim_pipe_pclk_in;               // DUT_pcie_tb:sim_pipe_pclk_in -> pcie_de_gen1_x8_ast128_inst:hip_pipe_sim_pipe_pclk_in
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_sim_pipe_rate;  // pcie_de_gen1_x8_ast128_inst:hip_pipe_sim_pipe_rate -> DUT_pcie_tb:sim_pipe_rate
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown3;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown3 -> DUT_pcie_tb:powerdown3
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown4;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown4 -> DUT_pcie_tb:powerdown4
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown5;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown5 -> DUT_pcie_tb:powerdown5
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown6;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown6 -> DUT_pcie_tb:powerdown6
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown0;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown0 -> DUT_pcie_tb:powerdown0
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown1;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown1 -> DUT_pcie_tb:powerdown1
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown2;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown2 -> DUT_pcie_tb:powerdown2
	wire         dut_pcie_tb_hip_pipe_rxvalid5;                       // DUT_pcie_tb:rxvalid5 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid5
	wire   [4:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_sim_ltssmstate; // pcie_de_gen1_x8_ast128_inst:hip_pipe_sim_ltssmstate -> DUT_pcie_tb:sim_ltssmstate
	wire         dut_pcie_tb_hip_pipe_rxvalid4;                       // DUT_pcie_tb:rxvalid4 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid4
	wire         dut_pcie_tb_hip_pipe_rxvalid3;                       // DUT_pcie_tb:rxvalid3 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid3
	wire         dut_pcie_tb_hip_pipe_rxvalid2;                       // DUT_pcie_tb:rxvalid2 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid2
	wire         dut_pcie_tb_hip_pipe_rxvalid1;                       // DUT_pcie_tb:rxvalid1 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid1
	wire         dut_pcie_tb_hip_pipe_rxvalid0;                       // DUT_pcie_tb:rxvalid0 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid0
	wire         dut_pcie_tb_hip_pipe_rxdatak2;                       // DUT_pcie_tb:rxdatak2 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak2
	wire         dut_pcie_tb_hip_pipe_rxdatak1;                       // DUT_pcie_tb:rxdatak1 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak1
	wire         dut_pcie_tb_hip_pipe_rxdatak0;                       // DUT_pcie_tb:rxdatak0 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak0
	wire         dut_pcie_tb_hip_pipe_rxdatak6;                       // DUT_pcie_tb:rxdatak6 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak6
	wire         dut_pcie_tb_hip_pipe_rxdatak5;                       // DUT_pcie_tb:rxdatak5 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak5
	wire         dut_pcie_tb_hip_pipe_rxdatak4;                       // DUT_pcie_tb:rxdatak4 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak4
	wire         dut_pcie_tb_hip_pipe_rxdatak3;                       // DUT_pcie_tb:rxdatak3 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak3
	wire   [1:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown7;     // pcie_de_gen1_x8_ast128_inst:hip_pipe_powerdown7 -> DUT_pcie_tb:powerdown7
	wire         dut_pcie_tb_hip_pipe_rxdatak7;                       // DUT_pcie_tb:rxdatak7 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdatak7
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus2;                      // DUT_pcie_tb:rxstatus2 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus2
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus3;                      // DUT_pcie_tb:rxstatus3 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus3
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus0;                      // DUT_pcie_tb:rxstatus0 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus0
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus1;                      // DUT_pcie_tb:rxstatus1 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus1
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus6;                      // DUT_pcie_tb:rxstatus6 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus6
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus7;                      // DUT_pcie_tb:rxstatus7 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus7
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus4;                      // DUT_pcie_tb:rxstatus4 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus4
	wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus5;                      // DUT_pcie_tb:rxstatus5 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxstatus5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing7;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing7 -> DUT_pcie_tb:txswing7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing6;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing6 -> DUT_pcie_tb:txswing6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing5;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing5 -> DUT_pcie_tb:txswing5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing4;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing4 -> DUT_pcie_tb:txswing4
	wire         dut_pcie_tb_hip_pipe_phystatus0;                     // DUT_pcie_tb:phystatus0 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus0
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing3;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing3 -> DUT_pcie_tb:txswing3
	wire         dut_pcie_tb_hip_pipe_phystatus1;                     // DUT_pcie_tb:phystatus1 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus1
	wire         dut_pcie_tb_hip_pipe_rxvalid7;                       // DUT_pcie_tb:rxvalid7 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing2;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing2 -> DUT_pcie_tb:txswing2
	wire         dut_pcie_tb_hip_pipe_phystatus2;                     // DUT_pcie_tb:phystatus2 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus2
	wire         dut_pcie_tb_hip_pipe_rxvalid6;                       // DUT_pcie_tb:rxvalid6 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxvalid6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing1;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing1 -> DUT_pcie_tb:txswing1
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing0;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txswing0 -> DUT_pcie_tb:txswing0
	wire         dut_pcie_tb_hip_pipe_phystatus3;                     // DUT_pcie_tb:phystatus3 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus3
	wire         dut_pcie_tb_hip_pipe_phystatus4;                     // DUT_pcie_tb:phystatus4 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus4
	wire         dut_pcie_tb_hip_pipe_phystatus5;                     // DUT_pcie_tb:phystatus5 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus5
	wire         dut_pcie_tb_hip_pipe_phystatus6;                     // DUT_pcie_tb:phystatus6 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus6
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel5; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel5 -> DUT_pcie_tb:eidleinfersel5
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin1;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin1 -> DUT_pcie_tb:txmargin1
	wire         dut_pcie_tb_hip_pipe_phystatus7;                     // DUT_pcie_tb:phystatus7 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_phystatus7
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel6; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel6 -> DUT_pcie_tb:eidleinfersel6
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin0;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin0 -> DUT_pcie_tb:txmargin0
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel7; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel7 -> DUT_pcie_tb:eidleinfersel7
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel1; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel1 -> DUT_pcie_tb:eidleinfersel1
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle5;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle5 -> DUT_pcie_tb:txelecidle5
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel2; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel2 -> DUT_pcie_tb:eidleinfersel2
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle6;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle6 -> DUT_pcie_tb:txelecidle6
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel3; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel3 -> DUT_pcie_tb:eidleinfersel3
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle7;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle7 -> DUT_pcie_tb:txelecidle7
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel4; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel4 -> DUT_pcie_tb:eidleinfersel4
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel0; // pcie_de_gen1_x8_ast128_inst:hip_pipe_eidleinfersel0 -> DUT_pcie_tb:eidleinfersel0
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata2;                        // DUT_pcie_tb:rxdata2 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata2
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata3;                        // DUT_pcie_tb:rxdata3 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata3
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata0;                        // DUT_pcie_tb:rxdata0 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata0
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle0;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle0 -> DUT_pcie_tb:txelecidle0
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata1;                        // DUT_pcie_tb:rxdata1 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata1
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle1;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle1 -> DUT_pcie_tb:txelecidle1
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata6;                        // DUT_pcie_tb:rxdata6 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle2;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle2 -> DUT_pcie_tb:txelecidle2
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata7;                        // DUT_pcie_tb:rxdata7 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle3;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle3 -> DUT_pcie_tb:txelecidle3
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata4;                        // DUT_pcie_tb:rxdata4 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata4
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle4;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txelecidle4 -> DUT_pcie_tb:txelecidle4
	wire   [7:0] dut_pcie_tb_hip_pipe_rxdata5;                        // DUT_pcie_tb:rxdata5 -> pcie_de_gen1_x8_ast128_inst:hip_pipe_rxdata5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx2;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx2 -> DUT_pcie_tb:txdetectrx2
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin5;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin5 -> DUT_pcie_tb:txmargin5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx1;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx1 -> DUT_pcie_tb:txdetectrx1
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin4;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin4 -> DUT_pcie_tb:txmargin4
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx4;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx4 -> DUT_pcie_tb:txdetectrx4
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin3;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin3 -> DUT_pcie_tb:txmargin3
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx3;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx3 -> DUT_pcie_tb:txdetectrx3
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin2;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin2 -> DUT_pcie_tb:txmargin2
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx0;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx0 -> DUT_pcie_tb:txdetectrx0
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin7;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin7 -> DUT_pcie_tb:txmargin7
	wire   [2:0] pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin6;      // pcie_de_gen1_x8_ast128_inst:hip_pipe_txmargin6 -> DUT_pcie_tb:txmargin6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx6;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx6 -> DUT_pcie_tb:txdetectrx6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx5;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx5 -> DUT_pcie_tb:txdetectrx5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx7;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdetectrx7 -> DUT_pcie_tb:txdetectrx7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak2;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak2 -> DUT_pcie_tb:txdatak2
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak1;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak1 -> DUT_pcie_tb:txdatak1
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak4;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak4 -> DUT_pcie_tb:txdatak4
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak3;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak3 -> DUT_pcie_tb:txdatak3
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity6;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity6 -> DUT_pcie_tb:rxpolarity6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak0;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak0 -> DUT_pcie_tb:txdatak0
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity7;    // pcie_de_gen1_x8_ast128_inst:hip_pipe_rxpolarity7 -> DUT_pcie_tb:rxpolarity7
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak6;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak6 -> DUT_pcie_tb:txdatak6
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak5;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak5 -> DUT_pcie_tb:txdatak5
	wire         pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak7;       // pcie_de_gen1_x8_ast128_inst:hip_pipe_txdatak7 -> DUT_pcie_tb:txdatak7
	wire         dut_pcie_tb_hip_serial_rx_in0;                       // DUT_pcie_tb:rx_in0 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in0
	wire         dut_pcie_tb_hip_serial_rx_in1;                       // DUT_pcie_tb:rx_in1 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in1
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out7;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out7 -> DUT_pcie_tb:tx_out7
	wire         dut_pcie_tb_hip_serial_rx_in2;                       // DUT_pcie_tb:rx_in2 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in2
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out6;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out6 -> DUT_pcie_tb:tx_out6
	wire         dut_pcie_tb_hip_serial_rx_in3;                       // DUT_pcie_tb:rx_in3 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in3
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out5;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out5 -> DUT_pcie_tb:tx_out5
	wire         dut_pcie_tb_hip_serial_rx_in4;                       // DUT_pcie_tb:rx_in4 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in4
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out4;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out4 -> DUT_pcie_tb:tx_out4
	wire         dut_pcie_tb_hip_serial_rx_in5;                       // DUT_pcie_tb:rx_in5 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in5
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out3;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out3 -> DUT_pcie_tb:tx_out3
	wire         dut_pcie_tb_hip_serial_rx_in6;                       // DUT_pcie_tb:rx_in6 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in6
	wire         dut_pcie_tb_hip_serial_rx_in7;                       // DUT_pcie_tb:rx_in7 -> pcie_de_gen1_x8_ast128_inst:hip_serial_rx_in7
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out2;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out2 -> DUT_pcie_tb:tx_out2
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out1;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out1 -> DUT_pcie_tb:tx_out1
	wire         pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out0;      // pcie_de_gen1_x8_ast128_inst:hip_serial_tx_out0 -> DUT_pcie_tb:tx_out0
	wire         dut_pcie_tb_npor_npor;                               // DUT_pcie_tb:npor -> pcie_de_gen1_x8_ast128_inst:pcie_rstn_npor
	wire         dut_pcie_tb_npor_pin_perst;                          // DUT_pcie_tb:pin_perst -> pcie_de_gen1_x8_ast128_inst:pcie_rstn_pin_perst
	wire         pcie_de_gen1_x8_ast128_inst_reset_bfm_reset_reset;   // pcie_de_gen1_x8_ast128_inst_reset_bfm:reset -> pcie_de_gen1_x8_ast128_inst:reset_reset_n

	altpcie_tbed_sv_hwtcl #(
		.lane_mask_hwtcl                      ("x8"),
		.gen123_lane_rate_mode_hwtcl          ("Gen1 (2.5 Gbps)"),
		.port_type_hwtcl                      ("Native endpoint"),
		.pll_refclk_freq_hwtcl                ("100 MHz"),
		.apps_type_hwtcl                      (2),
		.serial_sim_hwtcl                     (0),
		.enable_pipe32_sim_hwtcl              (0),
		.enable_tl_only_sim_hwtcl             (0),
		.deemphasis_enable_hwtcl              ("false"),
		.pld_clk_MHz                          (1250),
		.millisecond_cycle_count_hwtcl        (124250),
		.use_crc_forwarding_hwtcl             (0),
		.ecrc_check_capable_hwtcl             (0),
		.ecrc_gen_capable_hwtcl               (0),
		.enable_pipe32_phyip_ser_driver_hwtcl (0)
	) dut_pcie_tb (
		.npor             (dut_pcie_tb_npor_npor),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //       npor.npor
		.pin_perst        (dut_pcie_tb_npor_pin_perst),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //           .pin_perst
		.refclk           (dut_pcie_tb_refclk_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //     refclk.clk
		.sim_pipe_pclk_in (dut_pcie_tb_hip_pipe_sim_pipe_pclk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //   hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate    (pcie_de_gen1_x8_ast128_inst_hip_pipe_sim_pipe_rate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //           .sim_pipe_rate
		.sim_ltssmstate   (pcie_de_gen1_x8_ast128_inst_hip_pipe_sim_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .sim_ltssmstate
		.eidleinfersel0   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel0
		.eidleinfersel1   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel1
		.eidleinfersel2   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel2
		.eidleinfersel3   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel3
		.eidleinfersel4   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel4
		.eidleinfersel5   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel5
		.eidleinfersel6   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel6
		.eidleinfersel7   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .eidleinfersel7
		.powerdown0       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown0
		.powerdown1       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown1
		.powerdown2       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown2
		.powerdown3       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown3
		.powerdown4       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown4
		.powerdown5       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown5
		.powerdown6       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown6
		.powerdown7       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .powerdown7
		.rxpolarity0      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity0
		.rxpolarity1      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity1
		.rxpolarity2      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity2
		.rxpolarity3      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity3
		.rxpolarity4      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity4
		.rxpolarity5      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity5
		.rxpolarity6      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity6
		.rxpolarity7      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxpolarity7
		.txcompl0         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl0
		.txcompl1         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl1
		.txcompl2         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl2
		.txcompl3         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl3
		.txcompl4         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl4
		.txcompl5         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl5
		.txcompl6         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl6
		.txcompl7         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txcompl7
		.txdata0          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata0
		.txdata1          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata1
		.txdata2          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata2
		.txdata3          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata3
		.txdata4          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata4
		.txdata5          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata5
		.txdata6          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata6
		.txdata7          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .txdata7
		.txdatak0         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak0
		.txdatak1         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak1
		.txdatak2         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak2
		.txdatak3         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak3
		.txdatak4         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak4
		.txdatak5         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak5
		.txdatak6         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak6
		.txdatak7         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdatak7
		.txdetectrx0      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx0
		.txdetectrx1      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx1
		.txdetectrx2      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx2
		.txdetectrx3      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx3
		.txdetectrx4      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx4
		.txdetectrx5      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx5
		.txdetectrx6      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx6
		.txdetectrx7      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txdetectrx7
		.txelecidle0      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle0
		.txelecidle1      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle1
		.txelecidle2      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle2
		.txelecidle3      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle3
		.txelecidle4      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle4
		.txelecidle5      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle5
		.txelecidle6      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle6
		.txelecidle7      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .txelecidle7
		.txdeemph0        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph0
		.txdeemph1        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph1
		.txdeemph2        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph2
		.txdeemph3        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph3
		.txdeemph4        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph4
		.txdeemph5        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph5
		.txdeemph6        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph6
		.txdeemph7        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdeemph7
		.txmargin0        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin0
		.txmargin1        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin1
		.txmargin2        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin2
		.txmargin3        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin3
		.txmargin4        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin4
		.txmargin5        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin5
		.txmargin6        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin6
		.txmargin7        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txmargin7
		.txswing0         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing0
		.txswing1         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing1
		.txswing2         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing2
		.txswing3         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing3
		.txswing4         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing4
		.txswing5         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing5
		.txswing6         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing6
		.txswing7         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txswing7
		.phystatus0       (dut_pcie_tb_hip_pipe_phystatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus0
		.phystatus1       (dut_pcie_tb_hip_pipe_phystatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus1
		.phystatus2       (dut_pcie_tb_hip_pipe_phystatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus2
		.phystatus3       (dut_pcie_tb_hip_pipe_phystatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus3
		.phystatus4       (dut_pcie_tb_hip_pipe_phystatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus4
		.phystatus5       (dut_pcie_tb_hip_pipe_phystatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus5
		.phystatus6       (dut_pcie_tb_hip_pipe_phystatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus6
		.phystatus7       (dut_pcie_tb_hip_pipe_phystatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus7
		.rxdata0          (dut_pcie_tb_hip_pipe_rxdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata0
		.rxdata1          (dut_pcie_tb_hip_pipe_rxdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata1
		.rxdata2          (dut_pcie_tb_hip_pipe_rxdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata2
		.rxdata3          (dut_pcie_tb_hip_pipe_rxdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata3
		.rxdata4          (dut_pcie_tb_hip_pipe_rxdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata4
		.rxdata5          (dut_pcie_tb_hip_pipe_rxdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata5
		.rxdata6          (dut_pcie_tb_hip_pipe_rxdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata6
		.rxdata7          (dut_pcie_tb_hip_pipe_rxdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata7
		.rxdatak0         (dut_pcie_tb_hip_pipe_rxdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak0
		.rxdatak1         (dut_pcie_tb_hip_pipe_rxdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak1
		.rxdatak2         (dut_pcie_tb_hip_pipe_rxdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak2
		.rxdatak3         (dut_pcie_tb_hip_pipe_rxdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak3
		.rxdatak4         (dut_pcie_tb_hip_pipe_rxdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak4
		.rxdatak5         (dut_pcie_tb_hip_pipe_rxdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak5
		.rxdatak6         (dut_pcie_tb_hip_pipe_rxdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak6
		.rxdatak7         (dut_pcie_tb_hip_pipe_rxdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak7
		.rxelecidle0      (dut_pcie_tb_hip_pipe_rxelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle0
		.rxelecidle1      (dut_pcie_tb_hip_pipe_rxelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle1
		.rxelecidle2      (dut_pcie_tb_hip_pipe_rxelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle2
		.rxelecidle3      (dut_pcie_tb_hip_pipe_rxelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle3
		.rxelecidle4      (dut_pcie_tb_hip_pipe_rxelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle4
		.rxelecidle5      (dut_pcie_tb_hip_pipe_rxelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle5
		.rxelecidle6      (dut_pcie_tb_hip_pipe_rxelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle6
		.rxelecidle7      (dut_pcie_tb_hip_pipe_rxelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle7
		.rxstatus0        (dut_pcie_tb_hip_pipe_rxstatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus0
		.rxstatus1        (dut_pcie_tb_hip_pipe_rxstatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus1
		.rxstatus2        (dut_pcie_tb_hip_pipe_rxstatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus2
		.rxstatus3        (dut_pcie_tb_hip_pipe_rxstatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus3
		.rxstatus4        (dut_pcie_tb_hip_pipe_rxstatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus4
		.rxstatus5        (dut_pcie_tb_hip_pipe_rxstatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus5
		.rxstatus6        (dut_pcie_tb_hip_pipe_rxstatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus6
		.rxstatus7        (dut_pcie_tb_hip_pipe_rxstatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus7
		.rxvalid0         (dut_pcie_tb_hip_pipe_rxvalid0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid0
		.rxvalid1         (dut_pcie_tb_hip_pipe_rxvalid1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid1
		.rxvalid2         (dut_pcie_tb_hip_pipe_rxvalid2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid2
		.rxvalid3         (dut_pcie_tb_hip_pipe_rxvalid3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid3
		.rxvalid4         (dut_pcie_tb_hip_pipe_rxvalid4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid4
		.rxvalid5         (dut_pcie_tb_hip_pipe_rxvalid5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid5
		.rxvalid6         (dut_pcie_tb_hip_pipe_rxvalid6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid6
		.rxvalid7         (dut_pcie_tb_hip_pipe_rxvalid7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid7
		.rx_in0           (dut_pcie_tb_hip_serial_rx_in0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   // hip_serial.rx_in0
		.rx_in1           (dut_pcie_tb_hip_serial_rx_in1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rx_in1
		.rx_in2           (dut_pcie_tb_hip_serial_rx_in2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rx_in2
		.rx_in3           (dut_pcie_tb_hip_serial_rx_in3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rx_in3
		.rx_in4           (dut_pcie_tb_hip_serial_rx_in4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rx_in4
		.rx_in5           (dut_pcie_tb_hip_serial_rx_in5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rx_in5
		.rx_in6           (dut_pcie_tb_hip_serial_rx_in6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rx_in6
		.rx_in7           (dut_pcie_tb_hip_serial_rx_in7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rx_in7
		.tx_out0          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out0
		.tx_out1          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out1
		.tx_out2          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out2
		.tx_out3          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out3
		.tx_out4          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out4
		.tx_out5          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out5
		.tx_out6          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out6
		.tx_out7          (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .tx_out7
		.test_in          (dut_pcie_tb_hip_ctrl_test_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   hip_ctrl.test_in
		.simu_mode_pipe   (dut_pcie_tb_hip_ctrl_simu_mode_pipe),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .simu_mode_pipe
		.tlbfm_in         (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.tlbfm_out        ()                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 // (terminated)
	);

	pcie_de_gen1_x8_ast128 pcie_de_gen1_x8_ast128_inst (
		.clk_clk                   (pcie_de_gen1_x8_ast128_inst_clk_bfm_clk_clk),         //        clk.clk
		.hip_ctrl_test_in          (dut_pcie_tb_hip_ctrl_test_in),                        //   hip_ctrl.test_in
		.hip_ctrl_simu_mode_pipe   (dut_pcie_tb_hip_ctrl_simu_mode_pipe),                 //           .simu_mode_pipe
		.hip_pipe_sim_pipe_pclk_in (dut_pcie_tb_hip_pipe_sim_pipe_pclk_in),               //   hip_pipe.sim_pipe_pclk_in
		.hip_pipe_sim_pipe_rate    (pcie_de_gen1_x8_ast128_inst_hip_pipe_sim_pipe_rate),  //           .sim_pipe_rate
		.hip_pipe_sim_ltssmstate   (pcie_de_gen1_x8_ast128_inst_hip_pipe_sim_ltssmstate), //           .sim_ltssmstate
		.hip_pipe_eidleinfersel0   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel0), //           .eidleinfersel0
		.hip_pipe_eidleinfersel1   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel1), //           .eidleinfersel1
		.hip_pipe_eidleinfersel2   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel2), //           .eidleinfersel2
		.hip_pipe_eidleinfersel3   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel3), //           .eidleinfersel3
		.hip_pipe_eidleinfersel4   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel4), //           .eidleinfersel4
		.hip_pipe_eidleinfersel5   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel5), //           .eidleinfersel5
		.hip_pipe_eidleinfersel6   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel6), //           .eidleinfersel6
		.hip_pipe_eidleinfersel7   (pcie_de_gen1_x8_ast128_inst_hip_pipe_eidleinfersel7), //           .eidleinfersel7
		.hip_pipe_powerdown0       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown0),     //           .powerdown0
		.hip_pipe_powerdown1       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown1),     //           .powerdown1
		.hip_pipe_powerdown2       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown2),     //           .powerdown2
		.hip_pipe_powerdown3       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown3),     //           .powerdown3
		.hip_pipe_powerdown4       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown4),     //           .powerdown4
		.hip_pipe_powerdown5       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown5),     //           .powerdown5
		.hip_pipe_powerdown6       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown6),     //           .powerdown6
		.hip_pipe_powerdown7       (pcie_de_gen1_x8_ast128_inst_hip_pipe_powerdown7),     //           .powerdown7
		.hip_pipe_rxpolarity0      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity0),    //           .rxpolarity0
		.hip_pipe_rxpolarity1      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity1),    //           .rxpolarity1
		.hip_pipe_rxpolarity2      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity2),    //           .rxpolarity2
		.hip_pipe_rxpolarity3      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity3),    //           .rxpolarity3
		.hip_pipe_rxpolarity4      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity4),    //           .rxpolarity4
		.hip_pipe_rxpolarity5      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity5),    //           .rxpolarity5
		.hip_pipe_rxpolarity6      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity6),    //           .rxpolarity6
		.hip_pipe_rxpolarity7      (pcie_de_gen1_x8_ast128_inst_hip_pipe_rxpolarity7),    //           .rxpolarity7
		.hip_pipe_txcompl0         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl0),       //           .txcompl0
		.hip_pipe_txcompl1         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl1),       //           .txcompl1
		.hip_pipe_txcompl2         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl2),       //           .txcompl2
		.hip_pipe_txcompl3         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl3),       //           .txcompl3
		.hip_pipe_txcompl4         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl4),       //           .txcompl4
		.hip_pipe_txcompl5         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl5),       //           .txcompl5
		.hip_pipe_txcompl6         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl6),       //           .txcompl6
		.hip_pipe_txcompl7         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txcompl7),       //           .txcompl7
		.hip_pipe_txdata0          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata0),        //           .txdata0
		.hip_pipe_txdata1          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata1),        //           .txdata1
		.hip_pipe_txdata2          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata2),        //           .txdata2
		.hip_pipe_txdata3          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata3),        //           .txdata3
		.hip_pipe_txdata4          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata4),        //           .txdata4
		.hip_pipe_txdata5          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata5),        //           .txdata5
		.hip_pipe_txdata6          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata6),        //           .txdata6
		.hip_pipe_txdata7          (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdata7),        //           .txdata7
		.hip_pipe_txdatak0         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak0),       //           .txdatak0
		.hip_pipe_txdatak1         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak1),       //           .txdatak1
		.hip_pipe_txdatak2         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak2),       //           .txdatak2
		.hip_pipe_txdatak3         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak3),       //           .txdatak3
		.hip_pipe_txdatak4         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak4),       //           .txdatak4
		.hip_pipe_txdatak5         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak5),       //           .txdatak5
		.hip_pipe_txdatak6         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak6),       //           .txdatak6
		.hip_pipe_txdatak7         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdatak7),       //           .txdatak7
		.hip_pipe_txdetectrx0      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx0),    //           .txdetectrx0
		.hip_pipe_txdetectrx1      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx1),    //           .txdetectrx1
		.hip_pipe_txdetectrx2      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx2),    //           .txdetectrx2
		.hip_pipe_txdetectrx3      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx3),    //           .txdetectrx3
		.hip_pipe_txdetectrx4      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx4),    //           .txdetectrx4
		.hip_pipe_txdetectrx5      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx5),    //           .txdetectrx5
		.hip_pipe_txdetectrx6      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx6),    //           .txdetectrx6
		.hip_pipe_txdetectrx7      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdetectrx7),    //           .txdetectrx7
		.hip_pipe_txelecidle0      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle0),    //           .txelecidle0
		.hip_pipe_txelecidle1      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle1),    //           .txelecidle1
		.hip_pipe_txelecidle2      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle2),    //           .txelecidle2
		.hip_pipe_txelecidle3      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle3),    //           .txelecidle3
		.hip_pipe_txelecidle4      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle4),    //           .txelecidle4
		.hip_pipe_txelecidle5      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle5),    //           .txelecidle5
		.hip_pipe_txelecidle6      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle6),    //           .txelecidle6
		.hip_pipe_txelecidle7      (pcie_de_gen1_x8_ast128_inst_hip_pipe_txelecidle7),    //           .txelecidle7
		.hip_pipe_txdeemph0        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph0),      //           .txdeemph0
		.hip_pipe_txdeemph1        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph1),      //           .txdeemph1
		.hip_pipe_txdeemph2        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph2),      //           .txdeemph2
		.hip_pipe_txdeemph3        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph3),      //           .txdeemph3
		.hip_pipe_txdeemph4        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph4),      //           .txdeemph4
		.hip_pipe_txdeemph5        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph5),      //           .txdeemph5
		.hip_pipe_txdeemph6        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph6),      //           .txdeemph6
		.hip_pipe_txdeemph7        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txdeemph7),      //           .txdeemph7
		.hip_pipe_txmargin0        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin0),      //           .txmargin0
		.hip_pipe_txmargin1        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin1),      //           .txmargin1
		.hip_pipe_txmargin2        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin2),      //           .txmargin2
		.hip_pipe_txmargin3        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin3),      //           .txmargin3
		.hip_pipe_txmargin4        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin4),      //           .txmargin4
		.hip_pipe_txmargin5        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin5),      //           .txmargin5
		.hip_pipe_txmargin6        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin6),      //           .txmargin6
		.hip_pipe_txmargin7        (pcie_de_gen1_x8_ast128_inst_hip_pipe_txmargin7),      //           .txmargin7
		.hip_pipe_txswing0         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing0),       //           .txswing0
		.hip_pipe_txswing1         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing1),       //           .txswing1
		.hip_pipe_txswing2         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing2),       //           .txswing2
		.hip_pipe_txswing3         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing3),       //           .txswing3
		.hip_pipe_txswing4         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing4),       //           .txswing4
		.hip_pipe_txswing5         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing5),       //           .txswing5
		.hip_pipe_txswing6         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing6),       //           .txswing6
		.hip_pipe_txswing7         (pcie_de_gen1_x8_ast128_inst_hip_pipe_txswing7),       //           .txswing7
		.hip_pipe_phystatus0       (dut_pcie_tb_hip_pipe_phystatus0),                     //           .phystatus0
		.hip_pipe_phystatus1       (dut_pcie_tb_hip_pipe_phystatus1),                     //           .phystatus1
		.hip_pipe_phystatus2       (dut_pcie_tb_hip_pipe_phystatus2),                     //           .phystatus2
		.hip_pipe_phystatus3       (dut_pcie_tb_hip_pipe_phystatus3),                     //           .phystatus3
		.hip_pipe_phystatus4       (dut_pcie_tb_hip_pipe_phystatus4),                     //           .phystatus4
		.hip_pipe_phystatus5       (dut_pcie_tb_hip_pipe_phystatus5),                     //           .phystatus5
		.hip_pipe_phystatus6       (dut_pcie_tb_hip_pipe_phystatus6),                     //           .phystatus6
		.hip_pipe_phystatus7       (dut_pcie_tb_hip_pipe_phystatus7),                     //           .phystatus7
		.hip_pipe_rxdata0          (dut_pcie_tb_hip_pipe_rxdata0),                        //           .rxdata0
		.hip_pipe_rxdata1          (dut_pcie_tb_hip_pipe_rxdata1),                        //           .rxdata1
		.hip_pipe_rxdata2          (dut_pcie_tb_hip_pipe_rxdata2),                        //           .rxdata2
		.hip_pipe_rxdata3          (dut_pcie_tb_hip_pipe_rxdata3),                        //           .rxdata3
		.hip_pipe_rxdata4          (dut_pcie_tb_hip_pipe_rxdata4),                        //           .rxdata4
		.hip_pipe_rxdata5          (dut_pcie_tb_hip_pipe_rxdata5),                        //           .rxdata5
		.hip_pipe_rxdata6          (dut_pcie_tb_hip_pipe_rxdata6),                        //           .rxdata6
		.hip_pipe_rxdata7          (dut_pcie_tb_hip_pipe_rxdata7),                        //           .rxdata7
		.hip_pipe_rxdatak0         (dut_pcie_tb_hip_pipe_rxdatak0),                       //           .rxdatak0
		.hip_pipe_rxdatak1         (dut_pcie_tb_hip_pipe_rxdatak1),                       //           .rxdatak1
		.hip_pipe_rxdatak2         (dut_pcie_tb_hip_pipe_rxdatak2),                       //           .rxdatak2
		.hip_pipe_rxdatak3         (dut_pcie_tb_hip_pipe_rxdatak3),                       //           .rxdatak3
		.hip_pipe_rxdatak4         (dut_pcie_tb_hip_pipe_rxdatak4),                       //           .rxdatak4
		.hip_pipe_rxdatak5         (dut_pcie_tb_hip_pipe_rxdatak5),                       //           .rxdatak5
		.hip_pipe_rxdatak6         (dut_pcie_tb_hip_pipe_rxdatak6),                       //           .rxdatak6
		.hip_pipe_rxdatak7         (dut_pcie_tb_hip_pipe_rxdatak7),                       //           .rxdatak7
		.hip_pipe_rxelecidle0      (dut_pcie_tb_hip_pipe_rxelecidle0),                    //           .rxelecidle0
		.hip_pipe_rxelecidle1      (dut_pcie_tb_hip_pipe_rxelecidle1),                    //           .rxelecidle1
		.hip_pipe_rxelecidle2      (dut_pcie_tb_hip_pipe_rxelecidle2),                    //           .rxelecidle2
		.hip_pipe_rxelecidle3      (dut_pcie_tb_hip_pipe_rxelecidle3),                    //           .rxelecidle3
		.hip_pipe_rxelecidle4      (dut_pcie_tb_hip_pipe_rxelecidle4),                    //           .rxelecidle4
		.hip_pipe_rxelecidle5      (dut_pcie_tb_hip_pipe_rxelecidle5),                    //           .rxelecidle5
		.hip_pipe_rxelecidle6      (dut_pcie_tb_hip_pipe_rxelecidle6),                    //           .rxelecidle6
		.hip_pipe_rxelecidle7      (dut_pcie_tb_hip_pipe_rxelecidle7),                    //           .rxelecidle7
		.hip_pipe_rxstatus0        (dut_pcie_tb_hip_pipe_rxstatus0),                      //           .rxstatus0
		.hip_pipe_rxstatus1        (dut_pcie_tb_hip_pipe_rxstatus1),                      //           .rxstatus1
		.hip_pipe_rxstatus2        (dut_pcie_tb_hip_pipe_rxstatus2),                      //           .rxstatus2
		.hip_pipe_rxstatus3        (dut_pcie_tb_hip_pipe_rxstatus3),                      //           .rxstatus3
		.hip_pipe_rxstatus4        (dut_pcie_tb_hip_pipe_rxstatus4),                      //           .rxstatus4
		.hip_pipe_rxstatus5        (dut_pcie_tb_hip_pipe_rxstatus5),                      //           .rxstatus5
		.hip_pipe_rxstatus6        (dut_pcie_tb_hip_pipe_rxstatus6),                      //           .rxstatus6
		.hip_pipe_rxstatus7        (dut_pcie_tb_hip_pipe_rxstatus7),                      //           .rxstatus7
		.hip_pipe_rxvalid0         (dut_pcie_tb_hip_pipe_rxvalid0),                       //           .rxvalid0
		.hip_pipe_rxvalid1         (dut_pcie_tb_hip_pipe_rxvalid1),                       //           .rxvalid1
		.hip_pipe_rxvalid2         (dut_pcie_tb_hip_pipe_rxvalid2),                       //           .rxvalid2
		.hip_pipe_rxvalid3         (dut_pcie_tb_hip_pipe_rxvalid3),                       //           .rxvalid3
		.hip_pipe_rxvalid4         (dut_pcie_tb_hip_pipe_rxvalid4),                       //           .rxvalid4
		.hip_pipe_rxvalid5         (dut_pcie_tb_hip_pipe_rxvalid5),                       //           .rxvalid5
		.hip_pipe_rxvalid6         (dut_pcie_tb_hip_pipe_rxvalid6),                       //           .rxvalid6
		.hip_pipe_rxvalid7         (dut_pcie_tb_hip_pipe_rxvalid7),                       //           .rxvalid7
		.hip_serial_rx_in0         (dut_pcie_tb_hip_serial_rx_in0),                       // hip_serial.rx_in0
		.hip_serial_rx_in1         (dut_pcie_tb_hip_serial_rx_in1),                       //           .rx_in1
		.hip_serial_rx_in2         (dut_pcie_tb_hip_serial_rx_in2),                       //           .rx_in2
		.hip_serial_rx_in3         (dut_pcie_tb_hip_serial_rx_in3),                       //           .rx_in3
		.hip_serial_rx_in4         (dut_pcie_tb_hip_serial_rx_in4),                       //           .rx_in4
		.hip_serial_rx_in5         (dut_pcie_tb_hip_serial_rx_in5),                       //           .rx_in5
		.hip_serial_rx_in6         (dut_pcie_tb_hip_serial_rx_in6),                       //           .rx_in6
		.hip_serial_rx_in7         (dut_pcie_tb_hip_serial_rx_in7),                       //           .rx_in7
		.hip_serial_tx_out0        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out0),      //           .tx_out0
		.hip_serial_tx_out1        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out1),      //           .tx_out1
		.hip_serial_tx_out2        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out2),      //           .tx_out2
		.hip_serial_tx_out3        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out3),      //           .tx_out3
		.hip_serial_tx_out4        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out4),      //           .tx_out4
		.hip_serial_tx_out5        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out5),      //           .tx_out5
		.hip_serial_tx_out6        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out6),      //           .tx_out6
		.hip_serial_tx_out7        (pcie_de_gen1_x8_ast128_inst_hip_serial_tx_out7),      //           .tx_out7
		.pcie_rstn_npor            (dut_pcie_tb_npor_npor),                               //  pcie_rstn.npor
		.pcie_rstn_pin_perst       (dut_pcie_tb_npor_pin_perst),                          //           .pin_perst
		.refclk_clk                (dut_pcie_tb_refclk_clk),                              //     refclk.clk
		.reset_reset_n             (pcie_de_gen1_x8_ast128_inst_reset_bfm_reset_reset)    //      reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) pcie_de_gen1_x8_ast128_inst_clk_bfm (
		.clk (pcie_de_gen1_x8_ast128_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) pcie_de_gen1_x8_ast128_inst_reset_bfm (
		.reset (pcie_de_gen1_x8_ast128_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (pcie_de_gen1_x8_ast128_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
