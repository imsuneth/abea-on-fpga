// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:41 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iE1YOxWfka05EOly7kj8CrVAcpmRQJmQwVhX43vF1xXy1KHv+Hshe0V99et9SyG1
qLpVlTeMYcn/sdO0oBsCgWg9oJG1V5/oKGgE17NXYJsV8vZ5XigN/KkFqh8Urv6f
sMWEpiDMCJgv//lhYmumNiywQdFOHu28qHoa9JYX+Ik=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13168)
S8mBF4vVL2LYTbAVA4kAbTzZX2rObEcQBNWn57l6OLeaDlLdFTIjWJapsriBatJT
zoqc1kXof77sLeKkSQRU0KVVui2rqhYe4KcgOV8BivvqcL96jTvot0gqvZDgPYb6
kRgShZHZsiQGWxjKA1donTxXo3WREjg2lelNLP4wiVer6FWbGBLVj2V1Fn/igb5T
uKvG3TMMSAlkEI6rLNLfIu72xSkslQRviI+OVmy9eiudrmxirN8yYVvG1HaK8pFt
khCoXKVqvGSTkzRzC+5axsZEsC+IkmC/35NELuw0CvkL6lskC5vHr7gIxuF2m0yl
nraAhD4u2zagvMCxHPesw+tUZbTVpoRA8vNr1///Vhsj6XFBm3F7oa4yEp7WDpXL
buCWpc8/ugFfBiv8CeOss/SU5Qkf5DydkOXdYmHSSRdMwnHILjfI7yElKru7SGVo
24sYy4CfzPYc/kgTvIlSu8iVcoMGftja7ciSqgQ+wKXwA5EOEhkCKGFyLwyypMRG
ddaQgQXDY8YKKdlSeUzPFZx1ycqYXtBN/EjeF30iILHv7NNbEUkBqQxe0ztM5OF1
sjxmFk0jX08zoIDHNFhmtz0hN5aMgnWDQV98wf5FD3cNUBasNLDEBrXpOlgkUWN1
w/6xaBp/qZi4WFeUThHYE+qV1RGa617P7TbYX3RwQFtCzq388Z9qzFRCvLS1NZkT
mwMMGNEWhptXGYjxUNMaYe7YlT7ai8721AVrMBttPEuyMxk+wznFjeYMB8rQE4lF
BKMdFxueDJjRP0ZYjQtfU/0XIAqUj1unTx6YoYoKUOBiGcFM15wxBiOJxVI3wEui
DpNToBahJ+PQnOKa5U1WbGJqjaxTuA7+Jg4vxpXiYxu/QrTHGdxA0O/Tmf/jmQgt
8bdLUg1C58Ph3JBo8ZWT7SPikXacemGyf84OLQtKokzMRO6xf0LH5uzgeLYCY2Pl
IfCwd26MrFYdKNxcg33ac4RR3igotvKLSIcUocbILLTNvFAKt6ievydZyWddOk8W
qDqS+06ThsNQBSKe3Yb//uD4/dgFTAK8LRqwJZbIqbibSlOHkVdAaaLo/9JA/n5w
cYSaOtGSlhNMYE4aAZ1EzPS9wgjM4uhx3RSgcvY7FfVBoQN6RkaklkKn8JfWQZ6Q
fWuDPMZVnZHptXM7FhA5HV/ZzEvswp2utTGv7prrVXYfKp/9Jr/UVeMsVhY1UwpV
eKDiHCr87lQfEZrCRgdZ/Teq0sIWQtLtW0LubVidY1EyluOsuRSDMPWiPpJLrj7S
6xiq5GI50YhvFsoHNmQTqjZF7gkJtOMGnMecJSwv4FQNlEbTqmDEPvq3U5GKEJHo
8wHDVErPoBsVckvRZWXbbH/otUhfuDVi2PkWfc5eNOJ0g4EX0H8162gj7tvfmRR5
QDapmTX//WAr218ikMOXBDdOqU+rbsySlrgQg/+ZaJz3x9IEI+qIqCo4wHFPKwqR
zpnDYFPbjDCfJod4DiU/wpbr6iwHxSDbIOKCNy876RFgwiSAEQ6W2xD3WDtVB91j
XlKHfjjHNIQrosaDsdQ9HN/pvjD1G8SsfkfsZYufN2GY8a+fndHnhidKh098lJm6
f8bXEIZCoKvDXc8pI5WpilS3n1GNv+e9luX05iI452eup2vKBlix831sGXpLc20f
Tkr+d1yVjsWUDmsgCtkI9HxkII73eTjc1bK+eYUSeNLea1e8NAhR64tfXpXg80dK
zM3YFEMSYthXbX654Ls/LqwkS1Am/nLvSQLBlw7HmgAUbDx6suO6TM/T/Jb9T9Ti
ifq+R7vFfPZrhmdyqQM6WxxTKZCl1dVNNchFvyl/da10DaH7jhiAFZIzm1iFJwMH
Y2LhMzVUBhhBvEy6BT1JRM8pO2zj1n7rNVKkP5nEO248EXL7v7wDl+ftiZlgMN+h
4sgCx5iapIJSa2d2wOz3URgbJg0Omis4EPL+f+UzGI/K51cMM3aThIjRZVf/Isdm
y1/LtkOfPY0xyeYxyYF3CjTbWl+44sk71dIKTXrJWrvZ+qZf3AA4zn8+BtMw/sNc
lxpr5DG3SS28qZZm91Bfj+cV4jIKFUAx+XBQdRIZ3d/rIr7fCUjR3Sj8bmR7fkTp
vomDJJHtiUa8t9rWhh7oeKfTeikAMZd6zc80d84jDMZGjOXT8cezXkfuSPBCUeMb
vZehlhS5Jpo1rOWVTaOquWzXmX+gCoUPQqHjLCq/4P7Jr40AuhIzs8nFkoswV1JV
1ziX8t6TYJP0d5BnXQZsxo3TPD1RcJk+gdAhOXKU6GDTVkD3aXAToVozYIP1S980
+AjDBiEm8BeRrIaG8FOKqHobv4gvWX5ioPhHaSY8ZNWfhu8Qmh59lc3qPdynRTbq
KblhNtH/oJq1mcKtqpNft2X7SHXBsZFBZ8wgAa9X0qZ45/z/CyN928/EIvexsfLR
91vTXRwD1TVb0fvRLQiYvZRcPm9isCTKKRAWERjyzsa8pBmstD2VXK6AO47zB6Fn
SEeCsZgowAVV3uSadRummDPjFDXG7aP+IHxIl35EhhEpqil4cY1WIymrQr2fjNyr
J2zWi5zNtNEHC08w7J996OloWvTI2Qlq8NWgsNHzi2kAg/HtoR5Rx9Lg0nryrBjR
V4Rc9UmowjQzn+g38lLtrF9HpTKxW2k7mR6y+b1tAIIkL53iCPUVNgf/trdiNmrS
PjGAsyLXoA63+FnYb7iaIVQdTH3Bma6JZovGcKu6EPdsexAGMlRdnJpsAhjLJI2B
Zp9B7na6ow0U7u7C4bqLCRr84RgLEFBeW877PemIqIEv8a6mEYXSLyvqs8o1t7CT
sfsv/ucmg2K6Vprw3WH43Ae448XHIW4P6Hx2CHUO3Mhd8fTbig0QXVA+lZwBrO9P
CqaDO+YVf6kJ1ePEs4zry7NGXEBhol1BKXzm4GtqrQIpKZRehlzPtX74uBm/PEyz
OBYyjdz29mVJk1Z7HgKE90ktdrD3QAgmTzh0UQx5ahqOf31CRqXlKSTCAnpuuRbG
PKOKoycUG3Z96SvoI3Df6X0KJFylI6O7aLZivcz0SlMp86lODkS6SAJfsXqDDxXa
/53OIYjyssP8xYEQb+nxB32YGpWDcis/M52JKn47ySnKd1ea2BmdH3MVi5QxwlQl
Se7bJwt29AifGsWs8U/jYgmYzG11QOkosg4ckNiN3N5r58eowwnX0M0Z720CvRy2
oZNMzh0eR5OGmIwaRR3nj8ubhOoicj42zKeYvViNoMEWuUoCnwO3YBJo8+aeSyW5
c5qF1bxEdL8kcKngfVW1W8J5yzm/opmF3gP/jtOAQe3G1A052n/fL2GF9fRq+izr
YAxzqCzePguhl3hzok7xxfax7hjwol0Pye6aqI6KhFrYzU7GbaNGLIQjoAh3LO5x
iBIUmMn1ZwpS4UThb1MJEugZBuKm2qZrLMFa0TMt8IRjesZtnNMKQK2VY4goejqa
N0pnA9D58QWKnEoQjltpgvlGYIlcHYbF4X2pOoKYxxnUmR8UZYseXe0PpzYOYhML
qzE0EJzAmnqZsodHM3RFYdUcN3lefVyTdLBPDTB4vEoJi0w7ALrPUPmQMYQ83KWo
NAPfr1lzzbqfklKDqC+LiCjacAU8VquSgFPRXusIJ9YtSo709sfNc6RiM2eaQWok
IGsOHDqYyS9sAs/A7j9+Yvf2BZFmJMaBGYT5Z58NVdEEatRqbYR/7bDFpxHX7ApD
EmFKUbZ4Hcf5Kg2xpYgXL6YX/G15HICpFQFynil3VYHjQ530bRWubYwfR5DtY4/2
ViaEvW2ohBGsHHiZMsZgghUYbjRXPXszOt+QLzF6i9poVIm9lJr/I2mO6bL1K6Dz
5SiP3dAyUNc+smg9WBA3CzUj9EFUiwcyM1pSxUisGN9Qc3CsK9ak87pUJcnvlNHl
yhBfnCeXduSuN7QhsLv4/XHlKd3clWKJfBP65i+dMaq/GoHPuZHLkP7sdqUT0Ta2
rZI0Z8QwA2//LLhVQuqAhK+HKHytAR4RycoryObSXbNfppl/8u9pp2ahnkcfE07e
8hfQgf9dzmUfm87uhPbHKAtxCcRymjIM8XxT/JIUvIpD6BkKoFPOk3vHxXU8p64K
JNL1bM1R++nNgb0HCohqmQYdiGFUJhFs0/+NcPMzY/DmlMJNYx2jAhqikORjeGbw
gjb9JJrKjl9MDvu45QOwu4LDbpSIHzyuHTGCHQTEcM6Wa7IqvDHR+1T8fEUMxCoq
WdlDEEf8Eyj0RTcd/Vu8KAjvHGi+/5Zx71+qeujlcnn3s6/ow9xwVkVsP8P/EAVm
sIyAj/yW/kQO//dpuQ37K1zdY/DIzub/NWnLeNVec5iIrnR9gPtAktiXodqr8Yf1
oDqYKAidg4N3FDRXMDh5ovPlB2Phh87LGV41Xlm+cAI7ncOZvu4pTndjPRFWGWw3
b8YhHX7XJDKAr2WMQvBIUGJZRsvPPDFJvUX3nRlvvNvfRUdXYv8UWDPc6G1CvI+7
c0+93SU32wmJU+Y5Z6cxLE3Emu5T1X/+JOIkVNHU61JMVj/cO/XQWMBN49c8RBA+
4EdgYXa0Vb2gYrhlBnj9vdQFLurJ20MzPfVOOIK1Y6mvtpB0EhF8727nVHQ/ST1J
bDr63bEQ9ilAs6AsKpQu7K+9DRsLN+qCw7czvxedp2a2ckqWv3kn5ZQilZ9KoQD9
udlMIWnY+hF14osyD1lZ7FTgBfd38Qwv068Du6NymBia4GoFuTxhsjMBzDJ/RuS/
klcbGB9bBQg1p7ZaDgLlMt/wbea+4kni56kfcpZPB03XsZap54NyNd4gbLqEgXA4
4CcgXrWwcXBzK8WqKXcoWIMMGF61K0vZTWLgbRPSnzsYTBEH4eG2Sy+XevJ0sId5
myk3D8V4oUp3MoGsW0YYxd+z8erXPPV7t/a2fb0eyQWUoGOWKg5CGTGSG3jAUrZ9
im7/orN+d2UHLawgRxdqflsOBmsTk9Ofpm9Gl8jiQP4PFJdYheBgCbvstoFyFI9j
81TOjPXuRU6BLPK0oO7HoB+v+zCMia1JTjPjOnpIf0l2SGFXgiDryeGs8ipzt5Fm
410DE6MhVmJeMCPyxvTR35FOIAXUz70L8/G5mJvlRESx/Tf7MEGsxnzdOQy7mPg4
a+wUqphxsdRm1h2BSAS8veklHuMY80r9XvVjojOgPJs/RrICwbUG3BddEV4tHPQz
uMtd5KfrWnXBwPx2/slsKVt5tJK/TYq0aOU3/0lG3m6SSnYiaY8ZEWaKFNH8FNQo
GcpPN7jvCnC0gFEtgxW4k626QBZgPNMcl9QtBhaCwoHZ0OQT5JTLWthIJORosP5F
ZjFWfIUcS9d3O/LsPGVkT0GV9tZfHyUuG8RfyDd20fqfw4123FmwYHl7V4Qd4R+Y
kyiDcXWKqqZZMPPlb/Sfd8gnSe/8jXOi2WEuMHWBECCjVLeBD7BS+3R5EfM8jKbV
ABdrtTvDUaceXwC5tX3DSMk5JeevV7Gj0wC89bb5ka2a3An/rpNxf11/RSI4Bg8P
bjtl6HL8OZDkgrUSAgCcLeD+1IAy9mHfqK3WFmqcHnVq6PVNOEdWRYueyOBu7sUO
CK/EmQIjOKYf5GuPqfWqUe+TC152hhJAQjuyuq9pIB/XuY8gWW2wNuZLBYQ4AGwn
m2fvDDEGA3Qy6ZYnioWA9BZaIljUkUzxumrF6A6+qJu1AybfBe7jIRTxevamROxZ
BqZcqD5EoyZ156dID07IjG8FCZtyOBB8FlqFRKF7fa0IZJHEB1rndPFrB/lw8jRq
huCfzVqJl6L0RatkSMwkQC4nXHts1l4laWFQmaFlZ7iWVn4ntkEmFF8TPP0S0kv2
UxO0vL9frE7t/tEUYvnZfQZmIuufj2DnmuaLmZqJkEGf9TWljIGStmDsc8W43cux
lnAWj+d88nR1ssgvZ4T5HLgYkY0fVHkNSrTGCVAE3JJxtouW3CX6ZcIaM5gsNpxe
k2RthAxOFFHG8uTpeYUkLU9eQ12epDz6QL6MyomJUVoNjlYnj7U0P1KvyvhBg4ax
QpHEV3hxHpvKkoaD26otf6ZlSYpRDguLyXMQmCAu1ArcC+xqkO1aAWVVPCNV+oHZ
1k0L6qTzspUZQyQ+D8wOjE24d4w9lNpo8B1ALBZA/Cie090M9gMc8Vq4fgeVwjFL
+iqQKW3psDPMvpnv3G8Fk6xdawMH9MUyh/3RP2hCCq/zAPZwPZ5eBuEBMlYhThr+
SWntVUmKY+MZPcyCaWFYFGlJIHMJQceYnpL6Bqq4rZt0FTku5RCNN1Y+Ap/xYl34
gWByv+o4aG4DRW12ZX27AIIvjAC7CGGmth2ogFZKZnToAlR8YI4iGdtmgvTLuSVQ
20HvfWaOhiqXFnw9VCy9LWiRKwEJ6Fux9eQyFjAQberhxJK6XSmH8td33BpdsU2N
tfAckEmBSvMQBD4g0NCjSCrtZOv8MjqUUgItXTklL8xrwY4+xFifhAMNQG35fGF0
Q6oSoauGXAts3QwUIm3ffPmTMmLWEbynmPUH8pTT0V2K9PKZyvmRYeN6vj6I8t2V
n99zz31X8YOLlHoYdZRnA4chdJAPUsfuGpjvSYdf+x41b8wNboOL8C1v65p9mtwU
DAF0ThHXbxIqAuYrBYfQjgqCv8piIQHDdBlMaTUot9pvw3fBapCXQDTUzWWZG03u
mvJ3Qymkpc/83hYIxj6hIFV0OVDcTC2Dy0d24IGfhzIDNFjJldfG7kAYmaVuq6FS
t49rwEKCoua5asBn5JKeIQRE68UdQPUYiF23BwOTZrp8wZml2QJ5OfyKGtWl9k6q
S2wyA3PurON0+bk0jpDlyb+4Y/taDTmyiNj/9ZD+9I3gGqYHIEoaewY5nBLXEp0c
bV9XiXX8SLYCbAqzQBL2paHufHKUB2q4x8hCR9E1EUhOFC4UQvrDNz7wScr+ub6O
Mq3xYTvA+Az9xxGq/xkEhf0/mDV7zyLp/7mxwJFyY/LLsZtPcNWqogJXql7YvQDw
WS0QIJ42Sq+Kzg6kUcykJG80u2vCiPUSx/76PPEo5p/X3C9F4X3GUXiLqSpaW0L3
LSut0Qz8pWakIVWocn8f3tse1B9QTaYW5Kv64wPFjfvZwe+mtfqPLMu88RAO2Ka+
JHqpPZpU28RwFxoBUEAR3ODP4l6enPv6FMVTQMyy9lOGqdC6hBdBroMmoe3LTnXF
WMZbew+pfpsAXnfMHVv/+zvfU9Vsp/AUFK39rQh4nCp498Tyr3Gn6YwPkjvx4QHI
2qGtcR1Dge/r77GeTfCPxKFMUqt6x+iwEa0V7SpsWUsUZGJZ4KnUJhLkhAPAkbVd
yiQ3s3lvCO9Dndos2I9wjLDizHQRHhZYH1IDGem+HnwAbh9A+NPeAe5s34oNFUMA
YImw8zosZcieUJb3Aqy5w6EXCnAak7UlAlvHGvOovI7HUulbERBuJUOPp8Bk6nzj
XZXoZ2THUxlWsOrM1eLHryg2uL/yJimyr3g0VoKI0hH5T93EuMdj5+MwsJ/IwzQ2
AtxI/4iz7QhymXs6119/+yGGL/6p5m/iJKHzmMS+z59SzAYPzTX9OWrSeadyUr/x
V0Z6GO7xNIwZoGOyKQG574E46+3/BVbciwukaLhJ8tymO+VhsQfaydX0Hj9CFjf/
huAMX57wdzemxish+L1N4ZBviGWPF54f6geP4A2iKByGjevQFJZrvEulnxxATUPT
RQ1pCdAjqPjn1erUPV3EhZ+4EFNdG0Ula9WIMVG2uwWCujXQGLkxcmerscwTr/kn
Oh0i0FRmLNKaMXA23MqUiECru0oZWKmUvhoD90+9nCEYR+AH2Q8cCNVzbTSGhj2w
xVXqtmiAbEyIq2Wg0EODhbEhmlV+I5r1g9BTruIyl6vJLx2nANWx1NCyvxBOSnFA
KZDTcSpDR02x3P3WICXA9ZgE+sWrYZZ3WJoanzE2qMCTqr8z5DbBPG/wpyh2w1BB
dfx8J2j7dSWfspzfSmbkvU+LQDPHfEZJ4fc7e/9QqD1u3pn98HI0SB/9UOyXyfLL
nW7CaAc/rF9dEegOpvoPs1JAN89ECDTTcNbPN4zrjljhBljbD1tCqBg59VG3ar3V
3bYChdL2qNSwI/6M5qWsoCMCut8a5ZSEJAbC5eRBIorCsiULnkWr2LshAHxe0dL6
lTxL7hRMa4yfHHdrxWxeCm5QaBB0i4wldZtNNw9ozD3dBjWjh7HHB7irGX0lFsr5
qHbMkeItKFB1fTHDLithclfZjDaXMhek/EXJLUWj/MmOP6OhjOKuEZu13k3ZxlFA
RpvPrSFUw9idBVAr30V5h+QCB28xuzT10htawTjpjh4yz1o1QHSRpqPwj+JU3dLx
34gOMLMciN1/CsGMOFhKv/3O08MbJH0/j3HfhVjaqvfneF1LdNZiQ1GSd05NgfRq
RlLxRa5Y4tvSZF5OVE+hLFuXGLs6LtBhsWaT96SIBPZbAXxlzxgsAJt9LsZK2VUL
GI1xsciSBoTwrVzXwaCh0t5p3MyKwsYqqR0L4aH3D4yRfPNWIOFprtI25y3IGVh4
4XMyqdrbeTRoE7mSkYNEa5tqujZzVGyJOY1DtJquPpmIwULBP33+mw84yBfz6Np2
Vsr/SybgRfDK6UzhH6+vQNwX8wQU+XazEUvfcyfbq0e6KMMme1tIpYBJF8QbQIsx
czf9hvpofAj+X+0QagTSE2UgYabPrHUw5DPBadcfVdpuMHacz+1BWDszehuDEY0L
Vtxb+ep9rwy+EqpRq/YlVMJedSwa5mkm/+Z6ebdLXLP6KA8Xxzw82C65JamOauIW
ksVQydnAt4Jt6copISPVm+YDRUQhn7CWoVnbgp7svB2kft0JDlmZXfvyp1kYLtWl
EPtO55zR3oznxoL12Lfta0TXmmWA9592haSYCjYA0E9DZCVDs4wgBYrMjedj9BOp
zqGYM9krYPXc00WP35PPd94ubC5XbkU5bk68uE6JdQCkdn86IOHENhOtF6GDq0E3
BwDcGFJsOj91C58VJ1h3gnZpQaQmc4DesA7Ag4uHrcUkilJJ4KoP81PXiWj3Zrle
BQvSvNlTy3D+1J755DfExMmrqVRa08J26V3prCbSM1C3fjKkHN9q5VsOyH+ntUjw
S78dozqNqhLLeUetTQDJ3zPkf1AyoPeHwQtMNUtSqwU239MHBUiKq3dysMX8jTKX
IqWbq7Tc5WuXVdIYF02erjSuIbG90w34uJcVb/sUg+EP1K3xs809XbTIZtfoEWra
6XHVwr6e3UnDxkopQ4l1wzFX06j6xHs5DigcIBIRZRFI3vZ4v/bPiKSRCe5ToXYB
ubKpyjJkCg/8tezWpeIKivyqTwirpv40Jx9e2l5h22sG0t8n+jJDwumbyftmIsfb
B9bgKuzd+40++Y6iaP9q0KlezBRInHZYuYj7wE6fO/Ut9tmIivt+zT1x/9CGymtU
ERIdOz9DPdhVaAM1BxQPbF3P5KAo640ft0DSkyQYxAFiFDYgfPfBYPOfMUm7wdRs
DkBXiWQpa+FRlL8oygNrWAaqQ0i7f6MtVyF0p1KEjJJz07Dtu3e4iqM4nsXL878m
Wts/oU3aZAuEmp+v4dlbgrCI8lwbcWFQr/GJmEFAggqpFcbbC3RZuGMMYVgipmDl
lmslRrXsnOKis5eJll9YeeCf1y3u7Tgu5Lsr+vJcvr2i09J2RCC/0zzH/s/HhRgW
v1KVvYDsGP0RfUWoyGfo0K/Jpzn0seCKuB6jO0rtGA0NSMVMgdmE6EkDDut3gmuf
Qa+1wj4XRdhXfLzUt2nZIGfugBOciRyQj0TtEqK/M/xgrNxJE5+3EPyAuXl8KgVS
XK0tSn5Seuw7GCybzdH8jUAzOLOLIynpsac06xULK4Z+qkCSCPIKjNvVIMPD3t59
fRKxA1ASHs9lYlLXijxt8qi/ABayluRX6Ua2adeEV1pnDsww0uKfWc8wpuSUWJW1
Lpl1KmbzdiQIGL6eI51+mxSWXy+9YkA8G63TclaUROHbA8C6Vv5qPbt+t5JEDBh+
xEYuoDwNLWxERLMPRkEL/qwbmNJEEs9ICm2mdCnu0BCUud3/z3NUcYu4mBzRyFJR
pFIz7KKfAAmeVZeyB5ecEqonm4vYbIBFv8U615wi0aeQ7EuZIuw6/LppHpsPTQte
xIVymYsYbHiFPHMDIkiQgtHiKiziQU2YkHqfjUMKQG19w0LRLSldp9V81GwgTsFU
qCz29WCMxtqGJCtFYCe3oZeSUk1FLIxVAeW84M09O2tRmMaJOnpPmaDtbqvWZLpW
j6mBuWr1jUQpPHpiPz4qJ4nXQr1UbEIriAlZXUoaNfjJZl/4ikvdCWo0TtHg3dqq
6FAtfcy/iReddzOoDdMuKybUHf//xsKeZCCUD+EApQlgr7oeSZXggdGQ/FUbHxWE
EeHh4YxptTWam45DOM9rKMYe7US0zBWsVANwZfpQv3YE0nsUKH5nbSR+HjtBdw2f
FYkb0CL23fmWD0pb3lXU1SFd3CJFt475ge478lYp15etUt/hkotHIuCNJaN0ADRh
W/uOXpUFUAx02eCaxT1RzztwmUGPQDMP2ktZqgvzrGlxDFAuC9r++EzguMYz5xJ/
xZTHo2xuMxiWSkidt295m4ttQRntwWjyR428GMhlKeiWOePzFjWc0yzbmMlIoStx
29QdNGNV/CFBkdlTS+ElH8DjeIPRIoyq7gs6tw/iRfc+Kd7aMD5ywGcpYDCn45JH
TORoaea7YRiczW/zBQ7W0PY9ExLnnaviu1D3nn/lovolYYo3ZmP04ISZtzPECtQT
UxRaWuGQHQxBMGuquxZDDx5wAqAIixXH9kdg5nInscifk1egKFP8BCKX7PpmKW47
hu0mj8LXc+LA3C9WpEjBNrG1VuJBAn7AoAz32zh0W0GNDNMQTyFrsrp/POKU7JaS
kKBNe5N8QsLW009b27XcB3+/ZqsBGluiDkInT52EHBEKwb5Hlupf/z7VByaiOaWD
nfjpmdYCTSQbIb15de2MzEsylFgcn00Jxmpu6xazHUld56s70K7ODx91TgU6qPHL
m5Uqdnd1NSmsiuvVpZheVVnKFdBe4SaZ0A7kiffcggcykrtIIh4bRpv5joCoNoQe
DWFu/Y+3EWczfWDw6p1OCwSS0xpWGIWVTh5rxuCOP4u4giPbg9lv0pU4PLipUFzR
//uM18+u/U+4P/IN/U1ePDgFXVuVfXq7tEHoNFnOYp4fdMjQsR/6XuI5gnpnmL59
2vkDptkpHVbvnKqOfpHRgY/Lme4B5RmPOKnCtn4Ep7c/MDphmNfB3vZsJcQjemtf
VcbLxKz5grbvWug5nplJEvFviXcKLdGZHANr14UOf6HbXPHUjSsImDn4bky5kTOh
WnRjbVeoTDD2948uF7gdJnOuHcfvl6BV5wq/xrXvJOpr6cm/eWbythDjFiNFmR1+
UvOHFFYxaSOQivVxJX/mGenYBd61XkfU3+wh8mf9UU+CwQWhIGW/3kJGf6wH6uI1
5/qY3fdNAOJJ1gUHhP5OXQpQhCDW0o+zJKoNsNSyYLE/u6B3j3RncrhecQMlMTzp
fX5EwpbpuEPtCXg9kjAtk6elxNB6uwcimJqgWL55GkQsBNHpiXsrcm57mr1M6FvH
Cx9RZdGhr2gBQHY7ZLvQZM+IxsR/YHoQGEB9odkpcJW+iJKin52o7jQPCs4euD35
oJlIdHZqbYH8oJDP9yNnNz3sQf1d67+0+PzKV+40C8AkHkKRZfWhB/42lBsHh8zX
qs9NsyMYSjVOzTTuj9/PFomOTKhyXs5n6NWRR82S61GMEfShbEvjudL5He0ekX0Z
1Zejm2jIsJjzvvypifWXkhDlcxOAm7YSB4caoCtNYnOaIUUoSjxgxhfTr+L+ed91
WjwGtZiScijE44rRAQltCYiw+hZ1BCD8I3ypMKQN4QcpQ5mV7dCa5Z8MWQpI7CJ7
kuzsScTp9FY1fqYZagkyUj5WDQmGQRURDwVyK1owsMgcmWcYknmTsNyIdnolwH1b
UT5lVVR5ekFH37rLOq2oKkfQGWUYXI1idtKwhVbYC6IkDC9o7zjJg+UadpKpCT3Y
UhByx3AiV/6lORdNS+yjSb6aF9havHapB84V0AJUSGdW9//8mtUX//7upVMrvYCB
fhohSwwHpWubKjBO0l1SH1pE6BWO7d7K2hNZ+hSyFpwJAqNXq2ADDeEFgRC54KZw
jK3cZvJAkeVmmQ1CxyRsuTdrPyhJSqPm2uU5T1nMXKDzeUheyl+rMCGtWCZ2Jv0q
uheeK4ZuCjxT2C/grdie1LNcrrdbooFzN8XZpEPomRT19tuMwuclY5KnYkP2qa/Y
vjfNPyd7xrG8NPte6q5xWTJ6GoZM8wB8NDC5M7E4rKLrIBLNRMaEBORz/a8eZMke
TK43xVqA92aSlcCTnvVy9uOvYV7LHTdjoOemgpARNXqJdvRB6wESBQF7dzE5bybb
681qT9daocgX+298NiDaJjmQZi+9hV0NUoi/JwqlAFHiAvKo9vkCnCaeW6tEnrd0
pzSNodR2eSFXUUAJ0XQGuQalmP2lb0O1/Qut37/kfRgM7Q8hi1TxAw00frpyOmi1
0XWvLtF75yhidA+qoMYOm2qExiETrA/3nX76swR6uNUrFnwda6IwEH6EXtgaL/W9
/jAM1sylkzul5UiZH0MAQSVUk/Sn2HrrrClQAWV7mKuI4iraz2pPuZ+G931gXSzM
spqlDfY5qVuHMhog/cLllJ5rncFMpt0QaW6dcYRZSkrUAXFe+cRuXJutXN5SZTgX
EXxX34duKoDoEuVm1OrYx11x+2WyPTTV0y3LpS/pGlaa0v8J/ZvuPEcj8v62jcFf
+HhD5IMJvpnoxGFtCAG19tRBRaFZoL+E6vnUJRhhWk/Fu2tflXMOAhXePn9+Fi8s
kuihTc7v6IHhaj0+KUpUYQ5IQhvOueM6rmdXmUDEnZ8JRXNN8hrYnSbcWpIuGeXo
tFYbiiuGeSL1h9u0TeHyhDiaKToUG4f3nx3DAZtlpUVTDY7ixUJrI7zL2SOGT1xN
8+1cDIU/3dRPNtleKDFT2B7tW9e4FTy63oHdS+Z4Fjdvdk0FzwAEJKY2wcvXI6fq
q8Mx33+R10kdvakU7o44ZxIKk8PPlyHMTP2TDyIiYyIhMdnpCAuv2Fqmvuruoif+
Pw2Ow8l9CFDxWmvlc7fHdEQ4cIkX87uOYpSIoTtcijtEOJCKitkEpVkEOBmrY75n
W+kHSKYKmB3ka37qEuKK/OOpjuAD8RtRZoA1Py5IrwO0sP1nsv7vGMOCtw5ChnWN
+b58G61U071Fc77kFxtpjDXtOzNPYUHVBwnF7cRfEgTmjse9fJ4AlVVDsASj35kJ
hkWtEq+FRAxxKWGzjkJ+u0fEOcXe4bxj41Ftbln400IsGVlHDkH48TNSHW1LwsTT
qariwxlELqcaOrwQ2Ottt/vXmlZCME/sjF9e9xuI02e1vR3Qo8OXuqUuGK6RxnTs
vGkop8TChyH5vgj0xt6J0GidCM7+g5MoTtpwFHKueo6Vz7txUmfI1Fa232sPvKFa
9IDtL4wQ44ReIvvU8XXD+XsvzJYfQ7N5GMpuqkjtgJB974CVbE/Q016hj+lK7/3w
ytOs7Fhl6QkuZmk59ru1nghRhXk65U5qZ2gBXOsWPz3zI7Qqjdx8WQq2fSQQnWQn
aN1BbO+iNJSw8pguULBuLMC7v/gVJwhgqh+P9E9InpH3O8VZzrAjqMYwoG7fHnIm
fBFVwAaTwVSgTCJlcI+GgkK22aok4D2BSqXrNP7in3XlPw/vz4QcHmlOSkmxjtFi
riUlx+oyv9JXl9rxJHIYkMPENt1hNogxXqfHfxny8Q8dFGc9VmxxWmJNY/21l9Pm
Co0H5EZylBdDk1waDkg/8LHE4N5P71yNsqKj4RMFP6dimQvZF3V3jVfHkxElIcMV
paxCqPzMBSmjrgSfjBiAGwuIkJgiMV87Aqgu93D1pFFQrcKNl4sahfj5cfxxjiiI
nvL7Xe2PHoUIdbjxRByfedtTRhXDk/P8BKRFEY1SrsO/g8dmuFm1AatRRFsr351f
qwGjKEbE1mQA/Rbj7lPuVdqEvg46qV4/CGFBvC70QYiqpRXLUtNX4sqB0rrDqiqf
MffgwGHLVK3mpGuwHPzqfOFmNS5a21nNnc/TdQlqToafnaJ9lMION8P3GX+ZxGas
IR8LVzHruNjRtGYXUgGtv9gDiFIhjLGcPAiVDmm8PQZmW6uUtZhLSaheF8iSovBz
Uy+Xz73Rqc/L31+GN5U3GUCeVUQE96c3P5foNz/e76m3JbQhg1/OZC3EI8fhQbAw
dSUEp8kOKxqgMTYo4lo0Z7xcWfhBKoh0NNHb2Yybk+CsHMpkxQ3573eXNALUiukp
zQx0gPMZG92JwOwjyBBp9sXfhhTjKGtma1UpNl9yftBegHigDIfxkP56Vt9c8akk
jQ9+uc521mQ/M/qpY72FYuY3j0SV5q/Oph/BiAwiKtDaGZ0kkWAsbsmx0ucd2vom
YX1+2RLD6W0jqKCnvmiUTamuZYz/FI/blPMh+TslFmZbdJv5v8yMJONTb3qNH65+
ROinENJiGKZP1Ed2Lci9tm9RtOSpFH8dD3UindtuaLVeaRZcgOhTdlPlWvQWJ/mV
Og3bwiBKmFp2fHoEsCQJQM8r5ZYS1DYSVDby+3NOijbgA2sDIZBBeezMJLl1XvnJ
EmoDpuwtCXZSDy0JXOgCWh52G3hA69NgboiQ2dSaZoHG82Wq2sJRGYcmXDLYF+QV
b9ghAYaj4H6CYTvZITz1nlo3iHeBMl0iOThSSFezGzVsiaHJlNCZT/Rye+jINTS7
jK9G2bxJFzAOJ4Ipt7QsUTNMjLoiniFWuBbaEkrSCvz+t7ihbt8S3nK6lBzavdXM
T+hPYDZjJDRR/e6QEoIyZ+o9f8i8/7u+oqN4a1wK8Ao4ECvAX0Szgcm4fxEkUKyR
rSmfGo5yTz4jTds2zvXiK978qjmvbvMgVAYJSS5rPXwA1zs4GcKNQBbci3jJFbWs
sDUGaJrsa5Uz5pljlmunw4E4LT6nGM2mYFbmV26xxdeJv+lTDy01LzRCUGJd6axr
BpipLWEeKWVzMAyLsPKLXetLbTfa4pw+z/QyGYQ348l3JFGVY13iWrBLd0sk8OsB
DNECwaF+JoxsODv9Ki9doSWcWecI2tr4XWTPr5ySCAuYCaxyvmxcb0YGna5zzP+u
WP73cYonLJGHxCvLTFGrUYPP1bfpCFkXrwrbs4bfLmYqi99DBEfyRNL1NDBIZ3Xy
lTGKhO37Uyq5OW270Z3gfLw4U63gK38VL8iNrOPcstx2iSUTA9hktv1L5iFrqzT7
B/lKmc1bK3XTLXrJ/QpT6tfMzfptIdqFO6l2DC55xp4bi3Asrtp58nCwzzqELIbI
v4lW4FcllhjK1/P3xWbbxn2MjCF0+6hQkigYmh0Ar9yxJEcXBSB9j0QD/hbZ2Jqs
PZamQg4iULYgoTtQkfiys+Zf1AWWkdpd0QqsHah3u3ZK1zSESk5xGaZAlrI9UvHt
69UYcoLjDtWjAhq0WX5ItON2EtF31Xf2Fpz8knHJFULrb1dWPHTbXtjDtE/lUxs1
Gt4HSsSX0rR2WYmHL0pOIsMUiyejkf2tNTaM40xtucGcZwbczHWDxYWH7WW2J4OX
EdEQzrkVI37nbJW0fMw4E08UC+uK8W73Ds66UfriNMe7tdWSHxPRrAKeAe8b1HvJ
1h4qSbL0/MsqhnUqaLlIy9szJKL+VIDyiAY8zJ318/0kyomL5aETdje+GuErGjZX
RTmxcGiyTbPJu1KBAFCpT/kat7ca0etNZEthnrjQW3sCkS06QQluFi6Gex0E5AcD
8TYj+vR7dBnTDyfMaY6NFSI6Nbgi6kYVR8rYtKKYOyW9OMHDleIZ/xYB1o1bTuWi
RZXRifwuKUFrSBLoGyf+1mGeXPgo5SSfcWff2+vgJApsQ4V9mov9I+6CmYiQFq86
vEegv0yjTkuyR9guV6Z4Lr908A2c+KQYbkKQSTkzBvWtRF6NzhurnCvRyv10Y2UM
GmosAmYgmS7YCZAngGufr1947sk5PWO2zspCXkcXCfmIPLHRWExIsN/iOQEdons/
q0q65Q1x1/mWgOYi8PjBu27fa45hb7HPDIZM4EwMtpLCY1NOU0pCl6LFxNQTB4oE
hym4U7oUMhIVOHHgIuKih73o2JDLsyHN7C18b1LTvVo0yDlBjKrgxds8jG4P1L0C
ohHsN0ds0LCLCNPWjJs1LX69AmOjesRjUicaKAZbbEHuJQQKFIEiCadWSUZ/bjkB
flwqAdZ211WH4LdZpZfepDrl/0+0If+OR80c+FKHKXbf86Pym3yncssv1dKLj3Pb
ejN9zX8Dg2Omq4Re+SXr//qxeqd0lUq96bQH31ncZuvpS5WmDbLDcnad8DcPiBFq
kF/aj6zimTxd55R5Ji16B4MiGY3qwJLfXj72FeLicl7gxPOBKoGPh/RBCENYzJkX
ttp/CwwBmLlQVR1fvj0hv4R/1gfsypa4dObM9MDqP87L5Xqleo521FjBjSChjsBz
glnysWoXsjZrXk3c6PsU8+AzOcOhbCWTJXT68QNUC5kWBGFWBIXi/EHbs+wLHJyT
zEezi7A3IutEnoqQJCGhsTqe+XxGvUmmOCICgz5jcRKfllTbaHopNUl+3XQkHNZg
cs9EN4L5jToICxO2AtlxnjKL1619GZWuz5YRXmqAzSsY+jAPxCGWUJmOXUQqlHNG
salDWQIvrStZpAQGAj898QrXCgEP/Lwbma+e2XhKmF4zIs4q6+/PtIEnS6QmrN0C
+wJ6otRudghePw2nYGIZWRNOquiNrxkwo9arfHiutHfAwGTb9wLAWGW6FQSj+SUM
2tr85V59uLVmlBhfU+f6zmRe3dTyYJu0SOmVk0LPOByaHhZkOZQ3t4qQzg27RH7R
srkiJ7EKh8OgWUbmIMHsIXmipqN+sjc3XGO83Sm/lxu2nFf50fZpxJ2WRFEoyCIk
LYH2QXfYYboqysupjqNs3UULrjdRBepGptYQX+dQ/3HVsYHW7vbcCy4bQrWiADPw
t0K5rKqKPJ0ZJikJgRu60Im3RJPooFOfk/H0OVcCpb1kRYwcGyNor+QF/Nqz82Ti
Yy6zB/7e91ldqH3U/d0welIdKtIadIH95oer6LULTxdSi4VB4THRYaYB57dJSFMT
Vdc7Gh0+Bas5pXZAn55N/hJSWVeErPsZamZ6SPcLIrlIMrR8t3IHYI/QXf8clk/I
VyDIDzNIcAy9a/U423ZiCAjozXKW/z4PBXYnuq3tJqy6oj9O62vkJMxol+0eLMld
e8fx08B/prJpPiqbU5sZc45HneslM9Apgl5z6rpfErFHG7JIqaA1uSAonIrKcySo
xkDf5Y1QIXg5Hr62AZtGDfPvLGAmFitCsQnh+SsI3ZOsSHG5H9hPiS3uFkiDt6JC
FDyJx+WxP4134Gkg9wc0BcUysqJ2RzIW7JTzCiky1+1e9gmS+5xCha/GCcYFsieR
CDdkbhFj+islcdLVg6rVjwKTXSLHgfxm/nOiHbIO438tjnSpBLO/jDrrJqZXI9el
I/aNtDuzkU4QtvOgBFMIMw==
`pragma protect end_protected
