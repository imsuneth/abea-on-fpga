// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:03 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kSajno1Q0WAvCAVVC9qch9RVpgSZojQWQLr8/s8Q6tGH6c0mj6K0+i7PUZCOQ0JL
TGfuvJec3RF4ThAaqLtHpkCk8hQlY8c+qyXTcZWTEPTwjeTVmOErxS7zPc9W2m+L
tBsMCqcqXTnucG1iU6ZZDRa64oXt5Up15wS5T4C3/5I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
KzwJUS+bsXHQ6BTA5Q1dp/tEc3TcjWZQMpZLBz+21UCNFJU7Es5f7K82P8lat6zR
Cl9MzS/edLb3aLXFPTVfDYJBu1H4VZ6JSTmiZNBdK9ShggnibM7CF52Go5gDgDAu
6ue3b7omI44tQLz84Bm8sieBTq9j/hw3wVWc5iE068Zz+syP/xc+nFYZ5LqMyuQ8
W2sxDKW0St57zs9/Vqp6keMl2XunSJUSUXUVDfNQqtxQ4Rkig8nCwC968Ds9cIpq
2w9ihXbZUvhdfI0tVgS51tTYrfpBu9gijR6g0p6xCpHyghgRvyemAxRpA616/2wP
uMCKr14f183WDlUJ0anhNrjjBx5iYyNBSDby/SzaZaTgK4d20FxEOmUV3z/Vv1+N
9WMN3tYCYB/np4F9s/sKTDp4XqM2JzC+rynw5dymTgd4awOlCVOa+Mpns0ATubmg
8TnUiOR4MwORNvn+CcnHkLBGr1842qWXEkVg9SnT8eqXp814ySexgq3w6s1EG88/
Gg1CZCg2+NrkiJO/QaoGaJsP9K23YPuj/wOtZWj/GSa1AXk2w+7NjYGTnHU41PXK
K542tZIu7mHmgDqMCoN5YXdmDnkHRUqwJzxyNwY+UPPEsa1Qj0p2FXUdO1WN5hSV
Dxkk+ClYCBtuTu5s1nFBDqhHmJwkhWEI+fGrUhYQ+ctdJ3lTJNd/BC+g2ozMsPUA
5mahd9+0Q1cQeuzXJBXlFl9jvOToprZ2cWvyIPOWbzGhjkYlfB0Rfl5OGEz6wlno
UgAuK4QAxBbBfRJMl/9Es3EwsNN1FtVf1kAESzcnf2cmKkkwfwbDcXsAy/bCMnk0
yFM6WSjIEvTmCcd2n2ca7FI7f6ss/F2kkBRzMl8gaFEr/t6WAWEQULfVCHM1f7u2
RTPKYVAbGcyYJG+FiJf9JHsuR9YNAQN5O7GiYNdRMO96srud39xlFIrErvicSW7C
Ag4nlhdhVZwLGPWcWYK/vKH0DPzegI0CEeYLX1s6kc0ya07NYnqvZPv2BDOYjhDr
Y2q9DBgp8aA6hu4HTr0Rs5XWfVsFeTNe/OVel0MMIS8I7WMaCi12p45vYyGDJHJ4
q775JruyfjX8mawb3JTg7pBfM1mGa9/b3empVkbGbr4+FLPBCAb0PbUgzLNV/CQo
clPjiOSIiS16lxY4OYqy4xLyN2ZC2RrHt7rX4vZv3AeXvVH8aQc/77wX/TwLzVWh
M2+C8E+lgkHYaStH9USLxAJn5e92LPdOBbtiogWM4yExFsDcKOb8dzKgp0bhrL61
cIGbO+tAI8947vdPYtIQQ54bZV9SG+lnUeHYdX4aXkd+KEsrMS7PTqeTN4nRO6fI
WucCnOx0ysmygu34QlYlCfKbnSyVci4nNyC57mnsbMRQnX424aMGb6waY2r8irzZ
mMhBDm940JfINCPsxHeSURRX3yJd9GzMYyPJV8CNCL771SFuePIAno6H4SKSzlpG
EiQndKWwmDX26L9QtyNYD4wvkOgjmWUSOzvrEFIRKiVWplHYk3miDHpdFbYWTjD+
NsaiJjuVYseO+CQ0/fQJYS96+pDYF6+JjDDhDPsQCsTvAYH+kCyR02Uf0jB1HueB
Tm5FfF3P8SXGwn92Px8n8w2st5pyV1ltDQqUSBfSZdco6a9qfb5o5RotxURpLU6W
gDYYANg3rw6QG7SVbAtkfdwoyD9m9jIsw0Ribq3+UH/xJTTs2KnUNqyDIb//z8Rd
A/u7qQ6QogIRnwAMo12aKchD9rhEZsOsODNcwXQAcEmuKsPgn4sRhyJ9z+jUFPBS
YPhAlzhRMopnp7/cm/rHmJHLZOHFG0/+g1IKV34eakwe61ZK4FWPqr/g9iAJg5TM
Tzdt0cOHIEtx+0mkk3+oIy8SgFJUiTxfMGu62mdbR8HQko0TVi77yp+c33LEBbfI
Ygs+tTwW0NFqKShEThJoJ2R2gYiXNc7pcXwWusfZR25z3GwzfumcYqvAO2Ze2M3l
8A5ly8kQkzfczQ+LeS1zXhhoeTCj0dF/P7YS8WAjdum2WL1lbAURZcgpI3SPKTW4
vLHH23UPKWttVWR1+p4+X5gcNgeA64xjVMBnZQRd9xhyLUGPCfC7SeZCUbbK4dvw
MMfaYGqfdpEon05XHlbWUMmlbmP7gBStuWNrOzaqU403S8jZ/yV1NUyv9jXVbYmF
nQk7bm1RKC48YqKCFLMdm+3EWury8O02Myf7zXdKGamCrEkVA4OGarcnLD+mmzae
220DIOf8zjJlLJDzyDTDmOyVHXDvWO/qbXyYKwKz/iCRb6Aq4g5ldrRRqrCdrgR8
P/PJCE6anqiE4lFWTOpg7EJjO6RQpW7Vl66rE1P1+pdRj/nI45O0p4RrEaKAFh8Z
KUh9ska04r6PfKcmuuGmloJYbEQWqai2R4DjjGdgf4VX0FeqqG3j1f4w3beCcvUJ
8yC1fXjkgaQHDPw+MgIMuPsM0LmVeQUcgg6I0sYxVfV0u6p0r+2wQLM84Y1+0Gt6
+ATG3Z1ORJ5Y5GyX5z7HJ9FpzC5kP0hIOgQXEknCJsZpe7rGKGPSdRrjvkZ3MNbM
3P22gpKioXnw2PgigSQh5eP3KVmTJCUtdCK04PXRLREbHIPfM9awGDq5rSChsgPv
YGwSxWxjBbxkxw7fY3HG10DvTSuZFCDYwf30ZnQbl2Nz5sDkxXsxl2vuwRcxdEW1
BWb8xXdxu8KwMfg03yTERZGPu+OhVRlD2usaDyRPEDAZsPuRnCOz1eokGrWPC9lC
JX8hutqV51RTFNIQWgFmYA7UwzElbcERkAs8AGesCo6DT2wO/qz25sRmfxp6/v/J
pDlJvktGzsQHK8v+Cq4L+QwsJGJNfuPjijBnx3yG3jb3PcImb5fHVN451EYTYMeE
F4CTS2QpgSgiiZRnafL3Tt/rv/tZCYtDoD5Gx+0zHCWwbEqCLHexhkb6WGZJE71d
HOSTx8yoVFvD+A1ktgXlYPrsEc6H60Ih4JtPz61aTQExe2LgyrUMkH1btykqOLNn
1dUaN1KWaFDC+ZTs1QvWPv4m9onj6oc812Uge42UHTgeY215hlmL8tW1f8Nnms0u
nddrl7tCr4NGqVth2AD4/og2F55Ep+OKE6Jnf9CKf/iY/ny2WQrIrTewPHmabLVy
R9cDb+O8eK6m1JErCWBKm5Vr95sCJAU6V8MPFv4vurwts9RQh3In8FAl4yxijnpr
WeAZh2G5qSO7rqlZ/gL+5CSBD31oKDv0c1jFyaDOoWRYZwEtRGBqU/gQSN/D9utS
AXpdr/I6P4YWeilSE1/ZUhYWX+gVlSJ6yjUO0BxGzEHIx9bIYfyw6aNH46B9lomh
Tr3ykbvZsfXEIt+eznNhG1aYXfNqyzA86rbsFIbf9EkRTcLgKvCQ8OhIfS8kqHnx
uvI6zg3UaO8qubrdNSdqPbkgX5NFKENCepClJvyeJl6wk5/TwMOdtSh1A2ZFlhpe
jTUg0vYwDTgwvGUa26S4mXuAxxX2deQjEkepsf9h+WdqJ0zBNM4FGks6MnP9SVUq
m52gpUSICf7PVfPTWNKvqGfIh1Z3SztoziRrtj8faE5EAx3zDL5hQ5gVU8RM/+/F
oM/4xdOgmaiPyC95m8tIEQHip5ZlVoVQmu6rCasnHua3e22Y7svMm2hnNrXb5Z9q
cn89T9qDXAxY5uUe+mbT0Uwv47eFhNMIP7sIhM0eKdiO7CihcXSD6R52+d5/CX6q
PMFPN34ddhfNt++ebJJr0Y9mqXD4YQ+Uq+ZURtRGY2OFm2gUK2L5WciEytoD6Kw+
kpW+Kqa1f2/+0+1QcJl8DiqJe9bDI6xlY9ltmA7XR8m1qAs8ytlt43ibr0+Do/uE
w9Ft2TRuuULXgdTGe1R6Y5r/+3wfMB1mPd1uehS7Kf7+KiXU6zfWQ2rvz2pnpkON
YXzPB1M8QmucFKBdGW3wFo/YOYa3pRe8j9lTf+fbZCanNdhu8AjaPWTgR2rGEYCk
s0tL4q9liEaYJ6qO/FwpAIYTt76Ea3q109RuPQJ1nR1CNt81zopMf44q6zroqL7n
Wuws1o34n5kl1PiPEKvmq8Mi0/ZYr1iTDYzMkFNLxWCFIuWX87Ytxxq2o51X8eY3
v2x3FX/0c8OaofQIvy5l7VOJIiFERnMWOOAiobwmADUHOi+QHd59xSVnGX8K1vkL
WjSbe/TxNXCZucx/4EM6U4d2E6ljPXfdhEKJluvSZIcijYvKPJMwzLN4y7rCTS9n
Z+/0eNtxRjmyPd2J4gwUvB2QZiMw9/MnYJZhupAEDtgdH9nG4l1KSrrY2ggXchi2
aZU5gF7SEm4UHblz8rAA4UzO1zBcWSZhWySKvYzVfMsJf+vMw4n/UcOboB3hJTjW
lkk/xyj1+9asQq79LXLYlG9QMBsukvjmWqGckwxY+9aHf70b5RWJD+vR6hV9t9zv
jDGgOFOlvOJwDVoPdrxAEldULrIsPBzitR+bxxbliWdw0vmT3iaX26pB756SZnEo
t0ydguoZkdlzqzRrgpEUXGRXXQS89LSTDuy0V7XU//RcbrYWAA0Qvdgi7GGf4++e
8Vl8et/mHARy1N0RMVW1M9IA8ZvpLcOmSCyXu8ItUe88vIm+eh1rTMDX/UpiRMum
E8ugObGXadnpZWNXlL6zBRqs+mWovMy0fXVmwopP4cZwfi5oXiENg8l1qsDF9zO5
LNO+TDVtxl62kgHRp7ss5h49/sWDX5mVMuyuNAzOmJyk4gH1qWa8+uRHdg9SUjtV
qqXA81MGoz8HysubLcaJmsS2vjZAwJWBlc98UKiUUTlfqFabgPBKFhTINVzHU40e
RNl4Wf6zRZ7KUmgbwWXPQ5QW1tvin5M9qcjXAZ4UXfPAIEs9RQ3yTD953GOQ93yG
5Mpkqp83O40oWZ2w0/ttIMC1q/WhYt81surnZebjhk/OqUsqqPJSsoXodUFcUwOE
/R49XXmrHl/x+kSb1C6YyzqLuA1zNmWOtXm+MeSePDiTvXWPua+bLd/uFvWokg6A
obz4SbaldIKJJ6t6Z2CvnLoIEcFFHnnGEF3nZ9YeT2uNDERbUHrBcmpeTghkLH99
07ug8TxvR9sKVwDcjb79a3lbpVl0OmrlqQ9l8HdoNEJxDaJrVaMkpcz8TNUa/1UD
tvI0UQ2JoVqp/yWlZ2XP2Qai9CjQQPA7B8MKa6qKLOdfnrS7j7gAZ9VV1QOIoKk6
5EBQMME+d+Md2bSjWwtPgBKVx2rcyeTEjYs19ROWiy0h/ItZ6UvKo/sFD0VsXh91
xroEiL+GDSljHD8hfQLxOYWA0kmg26z/fxHyQoLMiRlCfWn+bm7YBqozdgZH2oII
bB8wyVuC4e+vgULwwe6IQU3S6WcIhLzGw6EP5FOwbBv3DreTiq3f/sEBhIbUnHDy
zg8eeeAN+nqrTEH2fzRBrYCMvqIYcMC+LlQ35a0vKSgtCRXKl1bIxFpL1r0wqL9o
z+6LebyL7DuqRFW251u96vqik1TQ7vByeB+WnvTxqJHtHlVP3nogJNI4SwzFE1bI
ftoRLLO5+/zloFQ07Lg4O8X+dyu5S9LS/ijVe5l7qgX29wlLjNlsx9GEcuey7lOW
rSfluadvtEy/B1gjDXoBc0ano8XFnTj0akUWDExbr2g3ksrmQJQwwW8r2xEdrj4A
ve2oQyTPY2lvAaO9+KATkAP66W88Au9rtA6xaDOrGCc2CRadh+G4XOP13cE690VK
wuHkIJGiQf4DD7OQJxmoJ2whej4WSOSKlXAyciObV49YnT9yJpdKMU/7vqpQ08ut
313aBYVfIHslLSJ1aGy4JA5iCPpyHWCLyXghjkJDVPAEBa834nWsX6sviSmn6HwX
ePBLFoJ+vMQr4oRXglxzHVX3tkWCn+sQhgdwdU3WZiTM/9Ddk29CC9cz1QAv+hru
Eio9yYLiqKDaurO7YuYM0TTwzBgJjwIMf5uCTw2lqD3IW0DwAh44nb5fyPXd1uvn
TkBghiUHLF51ctCCxSQbL+MMC34LEPxp4Mk+/vCxfa8blt1lg45hZWSyLWtnz8E6
IKi/R2oQoPYiaRn1OJ/7mcOC7XGuT59834vNtnsT9DJ+hCfZCENqBCmMgTSNik/h
q/JRdYKqDUdSEckRNlyndhW4CjygwTmbnw7KUAyem/F9CkdrSkQOy7aj2KVPBsZr
1Tn6HkUD0GuqlRhjeDz8lgAqBrl/VGtyhwzeBSS0jMk1mrPSznRAIfrfvmUPT3IF
WVWlum8mmSQ/K8GP09YjA0OzDummKqsZWVg+8jit0CQaG06wtNDSJKyX5hSUXT0X
DKNhL1VamN/S8yLWIQQW5o2w+4+Nw5dfXQjomE4c2s3DsnvB5cybkSeUPY6pybqk
jVs66BqtD/GEhQ0EYXgwIPsjnv7gxm7hytI7c6/eznEsKonG+5bGEGZ+ph9GaK59
if/N4kDdK1ONo2/A4RoRN7V5DvqxO3Ke+gYTNRAYL+glQyerCiNmcLAZPjdAunvn
2NJT+tsM84Fc8ZKNIM+sFzhacXy7amXvmFfw986/ZHdlVyYyxw4ZwnbE6QH6R+Vy
fh7WOZVJ7VTSABbrtgOCiBZgyn/FDguvgxVX8l4dT/v8pMslPwJZaO2jzMsxZ77z
78Jk2ixVdpD0tcR2QXx8UzVnA+1KcIXKxI7xSa3aPVSoYXEv1wHXtQln78uCL9fG
maWOcvQ5U16wUsqlLUKFSmDEL7aPO5Z2uTYodHr5AHX9L8UEFCrCfI/juKYo+Puq
x5Oi0cUSm6UOMiUkaY39DUdZcWA5c/+EXy6dlm0QJ850Y+KeumpR+nTWtTMnz/VY
oYDecrf79aNDR5958QKEV2rN9U84SS8Qrq5gYNmGVmzYqDid3WtGXJrNzP3ff4rH
G2JfBQWY/LDjJqNoNmZtJGowGyDpg1xhOfgJB+CPg3r+EHHD6C7/GghVEEbaIofw
QuX2eZ2xbKNp444sOLQYIzCGMXxv/3heOzEEPtcg9cbGGoGmEzW+4SNR9ittLASF
4WXnEDYEOXoKMFyW4NmF3UobZ5fSEIRzY8o8OR7azKcQfShcWZZWAgOuxa1igM/o
mQen5xJLqVLB9zHXLaBD+tyvAFsQdD5dy0FlktSZHHm574MbKfAi/RcIkX+WghLf
XJQhBn6DC5jux6SSvM+4Hc3LWe0e6jGaW3eN1OE0luCJ93hXC6FEmpHKI7bevwPh
WX4TqITG3JZkWEOvZtkhbOFDZNKVmswv+AfKbd5peztWgMqscm48f83SpxWXVblq
C90qHDNnKIAdy0A+qAK6E1b4S3B6sDshyF3fPmqt1PssewOu34/WgAZu8QKCqo8b
ogHRak/Rqx0WNcGRLgeQ9QTCDRn9gcsmZjzfcmxtjyCI0gbboSHWpLVLUsv4kBiD
0tUd3C1J4BF/5CIHmRocqZuEOwr5pHKLJg5DvImaQE/xYCYR0aUdtEvnsD/6Q0X9
GlEAjh5ktMaZLdGSNsa7dPMBKH1I5qnx2687IW23XzcuC6qKqjnwru9q+wWXi3dR
OOLy2zHwcl2YLgTa+z0ATE8p+msoS8tKS2mip29N48HPBGq75I2ugNhYzw6cIWbg
tDrgg+/oiz/TK9S5eoZZuwmGHa53OZ66PKBBT4tysf0bU3AbuC6bMQShJOZdlBZr
DJIi/cZCyTxTSRYoPCT2pT3uSRKrw9LSY0kssEEQOBW1nAHZGW/rhSHffch8NX6s
VZIdRLMftRho5gSz74OMFOw+JqGowSsQhBbor5IUt+G2NZMN+P7J7kV/iYl/CflG
pVxGhC65sGW8UzhtRp7AoddhS/63g81egmN0IP43L2bvdUV+ZAMj7Ao6FWghPM19
FkQp0wp6YWrdjBjb6OYBBT99gs6VmpOhOIOzlnwVbptnK0eM4/P497t++0gEmGiR
X7C5o1F3Khb6AmvC9L8qsnb2oyi6WUKQXFYJwJ1AvxFRu37UoQYfWPMGMOZ/FPC+
LznY7H8xgCNAP3GM+dPl78pxxUIx/+tsovYeDw9OCpCqMTNrTYoVhk7v0V5mDxC+
+qoyvpcEnNd1be5wRQ58THVznzEPUA50vXHlOful9jHnAl5TDgj+wrMcI2R3+yyQ
ZZjfoh2GJ9lz+A3798d4AJzKASj9J0U6CUVM8jij0B53nNqxVqqpFPxDGgU0JkYH
j1kqv6AZhb4n8YewGEa6pl63qnqYr6HLdSbO28KazPWmn06V8+nM1wCrRPv33XRl
w++Q/Vf+yXb4zcxWd0kTfA0o3GlB0JZEFbcYk7iqZAb6/eSVX6RBBOgzxGqBMR+5
sz1T1a/qOfIRezr//+WF/YCgxfmhekWAEwdpVEWx7Lg0lPR19XA4O/7fQR9p60sL
GAG5pBHp/ym0vzWhqehygeIgYmsZqxn95oVRZupuNCYAaiHjvRC0YO5PSdc+eNfl
6REWU+lQJWxVOZqK01Eta7f5csNaXUKWN1o2cm/uZdRXWZyf6MvwppXP/YxOk0Sn
NOQPBxiFuAV8LTx4MPu0iB8JftGEOcPLL4o6rDDDkGlvXO0len5n5Qdef706mfzG
gYvEOptG84JI5bewl9gsaA==
`pragma protect end_protected
