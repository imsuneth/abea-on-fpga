// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:41 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ix3CFKGIxHLPz1Wko5nrZT/+nzC7LLpHHn6qX2FzzbdsaohPEBVWkKq4263L4323
fx22SQIhaKkHdUpNLu9MfreiH8BXyr68PuVW7LC1QggHlYfM6elfyJQhiZMxLbDo
uCRWAHnrOsXviq/uIenwr+8XScJAIpF6EbtqUiCRLxc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2176)
vAWEqAFcm+vRo0cNXfQIBaYvGIo7i7VPr62uyxtBbFCNnjNVNt+JXKbeeDyfEdJ3
dSnCya4jt4YfMLopVlNAtpSVmAsSVLcT1ckCWcicA8quX3T21zaxmL/j4b0s8Ja2
9Lq1U22Eplt4QmKrauSFsRcKOsE+hBPlLXM5KYmJADMyJ1tE1yLvo1IpY4eBI0/W
EwCXFJnYkMOhFtRlUlviep2N6vBkdpvjFm9xi96eKbk5ontR1yvQfo7yQq1NStMM
MzrRh5nN3Tr4UkdtEf5dhu/EINFzRMaxXAFS/bPEnc6IHK5ARCQ7nfgVInSmUZ/g
eci4ciYrWbr7X5DWPjrCZZPPZQdrElf8L2m2ofx3gi4UTMol/078FDX2mGUGiUBB
E65ZYKofYTbLGg+C/jdLIbpJkVHTLwU1fmVE4gt3wXpfGzN9A4KvMx67FvzBLqk1
H8PIR7xQACBY7zO++hYwetJDOzR1zi+M5NTP0Rgr1XJAMCmUtaBuEEsRqyNaIiI7
RKjfLcivJ/JFkaapBz6PZ8HsRp7MnmBRZZv+EE7S0JmG3HJmGRalyQRoyE5wemVS
dm77Z8ayeFuUbDp9kySqN9ACo0JgBkVk0Y68LFDj+sCAkwOIkFntAKoZ0NjXDUbm
TMaSJQ+AK25d+enNDtJiowaEby1ZxNcfi2+cS7cWyTmr4qmonjDE+YyHSe++T0m7
oX/dFOzf05uuNiEoKUOp2L+JiDuM8qXUfYfdZwHAG5998vtqIUfscvafjZkb9mQ2
PoAwt3k9ZrZjKO+GqUDu7t/4N7daIwG6Nn/WPw/Sq/hnqU29chEGz4m5sv0ra2z+
FZz+U+t9cao+2bxxwVTDNm9BiDn9J4jg9+wGckqxaREdVOSaPq7GRUNoFxI7WfVo
ho2zkeopaSoIs9lPQGji5JI1E9awfsh6PjxHDyA+LOWr0dgzdg/dMMHZcGoUnU3R
bDxp/P+pW2sd8gw+c4ORdR56t2lhEvC95xIjo3xE3EstmdIEQgDMSkWlzpRLyHbV
xKF+WkBmeuH2mtt9nJENVli8iv53+FYG7eAFr7flZu8o0tGpnpwmtTf51qTXG0iz
o1TbfSo1JWEZBCVfNL2+zNFYQP16xP1C64fEiLXqvgVne/KK1FB7eU5KFlS34p/2
LsY6c1jelK0dhHGsF8AtKie3nLeIfGzCWSvx1XsyJbIJA/1OQ9ZtD0YBkIk2UVZn
FZTB6ikRUVVFVVhGOPodAAWrgAYzK/6lUl5ec/To2pEFB3jCB7PZI8W+US77hQtE
EDewj4/BgxPUJm4GPyHLK/N+/iuL4TXS4dPslFvmDYvLnUofWZLHHgQhFn7+XAqi
kr0eePTc/XZCIuNQHZ1DA2bqHfeI2MpSrfRVEYdVlgMMkn+CeS2t+HsV6axR+4RZ
OjzXQezBRzVpBXdGqwfPYaHXcdFDBvEB1kcJuNQgWYi9O5/NIR4klHqxOnz/QjYQ
Kb5jM+7svCu/4aU4abbqU8+swDqdaJfBdhQsovZO+mOgU9251GN+mb/vHOW0Ogya
95nglXyh6b/GC/XRuiT7shfgCuXNicuEKNnGLzaCpbu/cr+z6Y3aCrs4wxXHzbb9
vAaQKFzN3fMnHUen64+/DsoFxolfmaQGJAZwAZ+FpMGIJFThaJdDc6QKQec9E5mh
ZKxsZXysczxVZ8H+yyowdE9hHvp1oG3BGbzpOL1jbcRmaPRYlRvZiXA+oilAXrpn
vNf8Ber936od94CFKDIdzxa41ZMr7NcdGnkS2FpQlfJqXByyKqpQBb3pkeb5orma
HOoxD4e/OdVMgIRnPptOZ3X7QVhlZTrndvKm05rBA8wTLHcXKCeBCyEP5PBW/fxp
hUa6CxmOw8iP3imwWV0L3OuXsrL/qkVfPeZp1F2g9HkeGhYn7oQG4Zj4T0D1IBqf
UeyP3XmP4uZKKrE1zWrxOLnlpS5rmxykNZkDGBTnWFZRV8qvGdaQZCTmYQuIOvFM
0QDPZ1uHj7IlRISvOwR72WI6EyktNAdxFtR/Ci5G+ta+v4ZbIHriIMU/iENXEYqE
YfrRZ6YPXQV7kZCR4slc7gr4/EiY1lt5gLxSK+vKCn40G7SETz5ahgwlwhVgbaVd
6BC/EZryOdI+CGMnxtY3mCTlyp++URlAAidt4Yx01Sknxwwh3s+9bgxXJO1sGF/g
j91GwlWZ0P5L+vDONzzEUaTYPoYXyRZ3bySLgxhDMPXuEXEye8L5mUrMgO1XjuJh
8XhRIbYlUwnFbxSfzTAsPBg27woKdTA6Ztw+rWrF3c2jDUDXaI1aDct4r2C9AdW1
+TwK1/xb9h/6OlKKlPEx3FkCWDRQK3ed70FcHPNjGbQQuyi6LKyK7QTy4O4dsQTp
UDGrjy+gpea+VCib5MlGNqp9P66lCu394ZanV5HFyOEJUemPgMG1BfyFbIvF1N2/
QhSrbg0SMiK/DPd/BsSaGvXCPG1kh/lc92uqybJlKsBomd+wlbw9IA+xoSnajdMp
9N9KneufyLmVSDtDFgJfjDQ/YY4/pMLZrI9+mu7bupXIZ+ik8gTVXzjNF5BrZbjq
5BFG6fw+nJcA2eGPUYiWRxV3+S3msQbf7ZEpreZ4J8vMLo5wZOUb/tF2YkVP4hus
26j2SJoLMi3OzO6Rh+Cly2c6JtNaYIYjUl84hilIorAmckx8fIhBcRICgtmA2LWo
BIJqURH04kyK3RNU+pXa3ftEflGTD5FXjKsAr7rcar/IY2utRmsOJcIyXe9lSKte
X5osXEm8kWXxc1o/GspXv/ydECnbOATEvAkgkQ5kvoMWQ1ZfRK83H5Euog7dpCjt
6xHA8B7u3/oG+LvqLOU9dXEUBgLn7EHKnI+IfY2VlP6qJqSYMgNTu9D4AvpmjpI0
olxXCF5rAS+9/ZFKSqy81w==
`pragma protect end_protected
