// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:56 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GzQ4gRdEEkOjTHcHdjMjr+OrQroarg3llJlOJac02r0XcCmLvYy5yTM6ZnFiA8Sw
8OgPjhXYGBcvEpk8LT/PsKOqQiOBzRWRBrxWHFpA+kEH/aA9N3TvNJILxB67XiNq
QgUWVo7huH6x4BV2cTCLgW0T3minq16RucGcb4K1Eek=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3584)
abtNIExhUJz2ZNKQ/1J/oc+zdcafDsQ2q32fRBcwlRi3BTr979rfYi9uVQrQyFlP
S24laObd7cSf0vvZEINzatONMhuhmkZ8u5isQXxyCBzZNCHHPUFzqKm64sPvfxYy
9APc+Y3N/qfli6p9dYEnK/JEI8HEqpRABWs9OSiikaoqYgjva7BIlS6gW1yJ2sRW
I2UhTjw3ugof82WfILpOTqjxagn/KCiLaUGI/R6aeAO3XgkP/G+/4llTPc38LYPP
3RJjijdPcFcgWCR/1AdHBrZEBx5I4JivYx+fHo+PqewqIIU6lroG1OapbwWkqYS1
R0d9qPAq94wrCP9DySQYHMoH8fDU46q37vc9oNr7VJicmIpkntda1PfmHX4rr3dl
RcztJCxIAfSmaRWBp+v6dj15mFykeeL9NxJ8eDYsgkzbvZCq1YxbiaPJMwNPJg5f
mcQa6Ops19jS2ymoRQEs2tDX974BN+gSbfcE9ZBuPwgse74z4gpxMzJMNDDxh+5o
0TcdZtVCEGn6WgyaTx9wvEVRcN07yuO+NAZpx9VanHIVFj0TVBTlVtBmzdgmZ3V5
vMBbfrQYti9ZOWZ5/mtR0m9yrmD7JW6+HAt3EuHijvVGBEpBQewKd+qJwcYEwm0d
EJns8XWhBfMkAHuuvvV0vod6IGuTiEAO4nErg0DlFMaFPpaBlkVwET+FfbevTUDU
WxV/hAU7TfS452sbl1AndBvibl7xXZXLEulf2pyoRsR7C7C/E3HeVNoFHtSf/U27
HOw+QlRT9JiqKPOLYtqdjAar/x0zawQMUttb/3YbyVdTXnT0N4Y6Ck7HveFovqvq
8kN5x6TftjbkAM8Qa5FW9z6+v70Myugg47UwUBG9/K6numlnbcaSPfDJxXVZxXfo
pT8pX/6rk1Ab3nUONyejlS6DsteMqi/gjdw9AKZUeHZGXdIJFNDRbSow7E8R+dD2
1skAmI5eo+Ro29R5QnQdsnnhTzFf0JVt3ulmxAz6OTC/9duTdfe2tItTekp3W/xt
+70raolb/D/UYyYRqQG9ubeETfCXxdel4Ipu7XkVpi9ijAJd09ZfRFSMQI1fjYe6
vHlk92Y3TnXbVGjRvIE87d5Tc0cDvDvFPqlasTyxTkHoMbcTJCpFLe5ZebDe80b2
wHJWCWf99IGwawDtCGNSWhSDcbQxVKSscC+BbC9n4Jgp3VcFhEEysIp5w2w5H8Zq
QXg+7kr2y2DAelM4jvEb04YSbh+o66q9re1YALF2A5tszLp5lN2RI3uVv5au+LpP
ZeRrI348KbKgLVpy9b0vkrKme5a0M2p0f4BzgZ6Wjl9cdE3O/WnLm+SBIPysVQNe
qtQ4jafu3o1jJUppgPlpSKPYW7fzDk+8zSTELJUrSgwMQT23sfbyZiBNAVxXtH5m
zh/dyVYTIdrDQ+Vu7wpUhs7+Lk+7wvj1gg12tlAArqiflqqqtZeedeg0ZYlWW6Bc
i8dp59haZZtUXVusGFxusLBqgpUFZVRE9jqXpto3pyYsYGNbJBPUdpqfhSnxVvjj
SqZkicq6KmyiTxitpIzBB2oEUEzeLRtzj7oLzUkZdRuHc7hHS2F1yerGPyzL/c9n
6W+l06yJPggBH5d7BaIhOGPeOoZDGD+MGJ9349cIirgzz1kM/+xmSsCAp8aNgSab
K+sl3Ros9i8rB9si3N2A5csNgZY9N4PaY2o+TFg8Y7iX48NHmQsi6VhO1Mm43Ben
k49KCVE+icNEWxgoh3ivGwe5boe3AYlJtQQ0eRgGZhjMjRS6qdNYa8SwJvIztFZ7
B54K8CbxwOpdUpPjs+J8lju9lL+YqoHLr+qE3pYzNMbGePpDtJW0zuuDI8qEYUX0
UoD57Tm4yRPewpjJAJrajdEKpirFvcICeCcLVB9m1vh+RzwKVJMQRVsgSo3nz37g
pH5FPLBqfsuBOl2QugXC5Wso1lxLRlefXY9UGtHVxFljmmtHrvJnFH024hPumuYj
IZmsjbZevelTEhHLfApYGJV+ueZ/81Z6ILN/hrQeJQqzwFfCJqx9QGHCYnp2mK7Z
Is2hk62ezGt67ftKIuAQWThYY4K2lvvVfTR7lCJpjgOWooOOyIBeS5VqO8XAAKrE
VQxi7+T6wARry5OfFQQMP6cImsSTVooime/k5Ih2N0UBAHuUgC697gy1+Sq1murx
b7aG12MZkV1VOrSEqYsSDNdOHRXJ6/zxpJ8EqYvUqmrfLZNoJcNC0Xu+/PAkz165
/EancLByQ5Fvb3XX/Cj3nz3GIUU4PTR1+Uw5iJoT+B1fx3LYIfRKol7qDA4aH5Zj
LzROVlfivbO+oVoJa4aeypF47AH3nVnZff7a71MiMnXJ2ORKra7DkiQGTZSbXmuo
2wCX1+3lJWipHwRrFy8QnvVPMKx8czLz97galgaHi0FPWwzH6qCG012/VjqxZylh
SUBowCQvu7xy01lGAAhXM3xze3ZV5KsJS/y4WvIR7RR7DBfs+7DcPfEErEdSvF+X
4RTULyHlutdmLaoCm8M60pdaw2fuHAQOmelMbZBavqudLTGzPUCY6dPTFlTKwLz/
8JYzeqvkMnICZInxCXagi+xO3vQCU7+O/RjHjM6NfAWwr02vycWjGrj+pcv+C33+
HdjH32+k02ZK4LqJeAFmooeMuge4ATekEhB8yTkfLWbD9be5bOrcv8DqZZBN9Yep
7NDiHMVLZV55CDR4qMWVts87c2KRF5C4rugbr3RXzpoe1WHHE/lGcHMs9sXK2wtl
SjqjuhUnPJZqQUZvytvDA4UX0e4ykmOxhKVp4Gt6pZG9hdFvrHFG7g3YqxtrVVuC
F0DqaimU3qY/DWd9G8g56sMOCZDHPzCjAjJsFD/J/eyHgM7FaEk0k2w5AXUnxCLa
HuknzIVV8kHe2Move7MhweVNe5Xu+2aNGLBFaxBmjf/3T/+bFqZSo15z8TrnYp8k
RcdJBP+o41kMm48aSHudOMXt8sJRXt6IYQNd/tvJSXI4EQELlo4++Qc6OcwbjK8V
IH9JFsCUpMCvWA9aC8+5r3RzbeMBme9trqmVSUS7UZXLAqRTbhk8fXmg8Zpx/0DV
vRSyw4LDMOuI/lNn1JDwSaBsWriEnsN79car4TN0VXop7ieOX9QIxmgG8KcLXizv
j3B11VTYTtf7imna8yoNPs3MO2RUm1cGXVM2FacyQBx9MBJzdgzXhLzDGmHQe5yc
Vo4KG+DIKez7q/FZeZj2urosJ9MRTajCB33VoYgC+ibGs3WYyiNx1YJxoOTeVbOp
CiLXYWWGPyR8ezuei6bnVx+Sl3ulpizNG0n3iMYZC86t7tED10ZmJ9wjlDznumlr
vkfrdqdVn4TtOhTXJNl7/GbS7AtZAXC378k6QkBUf9nNgX6jb5jCSKluubIoZMbS
HuSDxZYYBT5DDq9PDjjCLt/geSH6xO2mWJcqfJsa4fUMC1EXHO9phXZJ5nCYygQK
MpGhKtRVh7AKJVdgF+fUhfbPZAdUJV2xmuit/r3lDQWzs2s2VCoEsLG/0KqNqgCK
Zyhj8QF+R452TqIywn5tCpa3+nNqGxDCblLUoxT9Bbg74KIeCVa+Yhj+/Fp5bOKV
PLAMIwav/lGy9OBN6WwPEHREm9N7RNSFLwrB40sU3pysK+dhuyNZqVK8iW06Ti/b
TJxAmi1Ub4AxOmedaLd+/rjvOGTaZbc5CLDqHAjpha6xmrPiAecyss+DVmszjeRZ
19rU1XW0eijDn8g7tupGwskrEmZRX3j9uVPUwEK/lnbtmLzT21pHJkC97VsfUaQm
30tMcANcdVEf9KCtbS9SR6yqIl7JNlO15ip4yBfZLcQpMm6prviJVE53mSm8nyPe
I5GprxOSyf/zADtRzMz3aSQN7ix+CCW4Xt60htPUTB7IG/D5/WhcFxwGbEnaYvy+
1Q7ajoHx5ZVGPpN1ebLNH9lX2UsXd+AkdtOjUZ6ZQj6VphgH6EAWo/70yMulmRAi
u6XewaFkmcxzK/hNhaKqKue/XS28ND702TRnZ0PGFvJ/43+oP5vBqsDjjAjOsNiL
oCidzOkahkMGzPoPSVwQlEzZ5pN81H/52rH3pA4yLasblv8dAYmjKvMwYaDwnqN4
DbzhdS8BDSJ6MJLNPRF6qp1xXLP30eh+RgqAShDu1ehbAzSESE2VRVp0ZOZAKayM
bZuhACHG3C4nlaZCt/wGIh60Yk7LIunsenX74qmoT2eZsFRke2iEf0muSJ4tJ3ys
OJCUqE7/V/Mhv793FA3iqVZLhFKALwjTISKMSFU336i5IrkC55jcy5ihTeHQ42lB
qwP3EfQlCWgoeDFaJjjxZAdTGZNHPwIro40zaTA+bJbGOjcT5QOTuGicDjzupFmd
b0lX3K8eANlpcBVmQqn3jWLSmMoRCKNkN966JTZXt1v17y1T4zTJG2pHkW+uvGZ9
NE3l0XwTzkstiauKBX269L9LwAlcTef8XqNGJy5ECSc79pMTiimgmblQKAxyHGJL
gearDvDcTACStcNRH7t1Dmcn9lUb20S9Fmbta2X8y1N9VkIHtkjMiE5wJWLlnzV2
JeJzKHB8jWY3sfYN+kZ+TDPTX666qOLHmoGs6OnTx2uyWHya1gTLZmySNIeuAQt8
baFSpMVyCRb+ZH69RBQMPw4qDH2+qeRNnb2v8/8xhj7xqZRBizxC8Z+2PQ8kBrPq
/YRl1JdQwI5WpCq+cW6KRhF60u++PKi5w1TPlrKThUbPjJdrtZeJQC2PJtKHOR1u
+YMbn1d8MYawOdFdk8f+rQsyQYbk3pEr33F+4QLfSRc=
`pragma protect end_protected
