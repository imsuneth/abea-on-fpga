// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:31 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HMZkgMGkCcfQchXn039cE+skjAMwT1KQbOnUEaxE76HNyyqS84jQox9PlDdFC1Bw
2DbXiekWKavet4zLhYRVwXzUOSKutCpA56a/AGL+gbPUGNJin/qsH7DY3OgBHbDN
pdzw27sMmrEBstTpTg+h4zKBiDRcKnpnZYFfC2abyHk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5552)
dB2xCAJPkPKKvmhOX3HOd1KrPajg/MOly2ZYY/aslIbMg/X/6W23a/VU4tUG7HOX
PzY9H5S7J4IVq3wMHccMnlcOUFAGrYzErMu3q7CW/h+S/9+Y1O3GfLlKZWYXENvB
AojEh0xpYNC/T3xCVlGnSNlHsTA9LOIP1q2b1VnuNWw1NP0/sx6odLKlooEoeBcm
JpoPoiJ94ZMCEGgGmTSod/JBAOrddCQur0e4RoxNZBrBO6ydgxJW9FqtGEvtfzKN
xJ+t0kZ0tgp0I9tYDb4La/+t2Y5//ogzXvx0Tq6vf+S7asMz5Ujet11cXnmKhjFx
gt/VkF5kpysKjFkGGHqCl5C9hYRVmu2gkPNLeC0HWcjjU77jXL8WQJSyLOEashPx
f+MwH2VEHqNMnUmilstGXnIngfYhe0IhsoPTwbArbj1JNAeQxv9x/hmXXOQdSFky
Fzk4KLHgGggpOpGz3wlEe+UsYuiw3YSLtt0AdQ8esU9KhxY4NTX4x23gMqCv95Eh
irt6tozGdJ0F1Q7N54triEhWE+G+ES5/lsgfURA0sJ9vIlxZb5EC/7aZrgJ44fhf
vs9iYqIXGMLj8ppwgMYWlXBRO2YAn2AMCtrDy7/iIiQrydRX8umLXWs62HTRFyhC
307NT1Tw0KU82pTX/dMupiUu+21gPMpZbZoTgqPhxt6aRRdLj1dUTDYgrs2pkARg
EgCsbzFj+q8S1emrlY/BRMh7Pm9+aBNFUHODdz/KqStwhSR8lJJmNY0Vrbv0HFrx
A58Gnj52qcKgsGPBhb6FlkuyyofqrPG1HY3vBq1XBti+yeKEZFTpLdS2YlHS7MQo
uJcT6dpKn7T5IONoZHtifLYJ5l1GnGmkjDQ0y1ufQ0KroNMz9fBDEaqLHrNYA5nC
eoQXDlZ0Nz2Uw1ngmiy/EsCHFbHnSWxR6UPW0ykEuj7WEe2SogVezrcSr3h9ymIk
7UVD3gtZMEiAzX41YQXDd2+XnN0cWwW28nIxODgcIlcLRiH/I61PIousYDKPL7IO
ayEg5VD5Pq8xbWLsGdiifzZQtfShcAreAheDaLsTkOhp6BvI4dlg6wiDvPWKaf1F
OviscdbkXkHABYio2eb9+QDjtFBJCKmMsrbsQyfhQ9fCEHO6Hi7wt1wPRwPZ6nHh
gETCw+xqFoMVtppEMkQuoF3n0cocLaVWdBUE2/KdjFBa90ZuWig4oz7naHHuSldp
tEgNFYK5+zoVpoaMSO4Ky9eogSQOAp4PB5El28lX9+3zeHrsCpIq2W5oxvQXc1EV
kAacwsXIV7lm++enIgzR17S1VIWuScLP2R3xZMRMGRkhXvgbvrqoc5AS1geU/tdm
gpQyynF18pxdMplp06+Hebgwc8j39/dhcqUXs62TC908I1Mho+Nd69VxmFtVXQUI
of2phV5uASSwO0u8ckmTG+h4L9H9sIIgm0dOLC2iaeMSxL9K6c6Ifw5ieETZew7q
x4QyazcIZvGnNtlc2OYA5LkEcHb+rmaFu5Hjn8R+sP0/eQwgHtM1XyRqcr2cA4Lv
KcO3uKBdSrxpVs1vNERrbvyv6poOaghtE7l5kh8rxczYJAo2+RtuEvQTyLuFDHCU
hyoNesDxZYKvZRl7ATXpIrJB2wcUVFATXorh6MQh5qHuN5NkxzPV8bEtF/2GlC+P
G8efofJUn5Q6r+NYmxWsVzR83uzHAw4b7qjzPdXLHbBGSIgnovSrToKYgUnfDj4j
nH1CGAqPIYEkdPIKsJSp+kbRScsxDGvmjqnHicFcazespsMyRmYi41T6Ac3h7FKe
PesKMWaQFuCsXPQylqIVwATLYYAM70EywCYL9BawBb5C32a0oTr7mIYvxzrI5+uh
3yc10Hy4A9EVnc4TLQ/NaqLTJF7UsqcRUoREVlVFfGbpwY9eyKxmx4UA9v+OTOva
z6SZyn+LsEXEekzZ98kDPH0xRNLfk2M7HYM3qASxe7BJMs5OxCbYZo7uWT+tgQRW
I5lQ0aSE9ZNbrT6AYx0D189iGumTFncgJCVSQ9o1QTLkaosPIc6XBc7j1cp2S1mQ
wQN023XgI8cL58QKzIqAQMjNtmNnbDWg+RFEuBhtPnJkzNm3htaosjr9LWbu3r9X
ab4HgKyPerAQ2YE0y7QhIO6YwZwutOJ84o93IXbHkGYI6x9UKuCLUcKIFcxNy3vI
NFqIF/2iSED1Zr3BIy9HwcmcYTZXZwmIPArWvuk2XIgWR1vf52mJ28Irqb+X6LdQ
aLVfwWCeSLD7P8ZHqONCUEKaw93AcuTU6YY16B1zEcWH9hNz3g4RV66gbkH7F2xk
KPM5OjQSIbOc1JyKvzig4eFSF4wOZfT8NZisl374TDjzyNTsW6RZtiqA3kFUQT8q
TqKIEKvatrP++R4W7aDptmZ5f3jgMd00bflmG+xYi2hfEm60hHDv3o1C1rROMh5I
t0qzw8MfAdwS0mHszbK3fo2m4mOIFbW9Pu4x3PgFNA4ufwHW7rahL2dA+2rkSIc6
jUVhIUXtG7WrZrtDi9+s1rqO29PR2LysuQY5gHJzMU/nJyK75AzxpBFB7dJ3jBks
d0Y2YmFM1pyMY2J+o/ETo6QpkGtczdlr8lZ1AcnXfCBg0hRJXSvqRYdZIX5iruYb
crgPN235jZ6f8F9qRDfOP5Wrsk4aHjMMjcYIB/PnRoAZtqWbDpgQt0S/UzHU8B+e
bRHrBl0wLRe+Loq1+uMqlEH1ZwRCka+FiP5LSqHv6n5u8ZZ7Rm8ApSxSrdZ0G/wf
US53DSxKGgfscnli58MBahM33+g55WVT2SKR7CaWzF9SIHHvsO3ZtMLZYxIKSvh4
ZbMGjbHRdAg+a+QHg2AzAn60W8bpXrN767YnJvlHPBZjP2TwYi+C39vmfjT6et6T
z9xK/K6I8mLzEt5sk7VEz4imfdyW7J7vqIz6umsSmHyFt4U/jEj914IKJQm5gtQE
MzRxqIUvxs24rQ5kDgQeAmkIfLZ71oKSQ11lOVVoEyVLtmdBPF/a3z8J6E/zS6il
9WAC6UcA0Q9s+v5YpynfcMyN58LoC17kvYvu93udJ2fH7vLIxHEeKJ4ic9w4TPAp
FueLyk/fWOc/tkeRJyV9FfT3Rn6DZiLnq4LDmlJaooHYeR6BNq5Feo5RajzI6iV3
NJBESynyZH6F4hxItjWqy/1eG6hq2ttKcD/KhNyZs5ydG75EmD3RyhA3wHvoN9A5
OPp6ZkC3xQcwCNF4T8EH2NFtjLKDJzSQUolQUSYPcvhH4OyfSTOmc/94xx+/h2mb
Me8KYx8V0qzVogkjhmk/yRyK3S17WHx7nZ0dvckrW1y80+N3e7zcTwthbp9EiGG5
QB+kJksvcUL0/NN4c0Dmdgeqe6oyC0HcvxwlWuDbAJn31FXCGNYWROMQrf4w0boJ
hum8TAO669MGU+jrZUg79CbvShvk1l4d8UVCztkQ7j5aISlOlDE/sDbD3e6cQwvs
eAqNeKglNvYKW708tSgypliswkqbCJDkWxwDDFGseffbYJrUHeQAFPC85dSfaRkU
R6dO0FC7q93xOnmIKAu84ZnOZsx2hG1Kg4mbQH+TYGNUXmn7SyvLYIqR9pSUTJnj
fmtPjF3cAoWytWW4tEWgjrPOZMUABzpVM8Ae2jjZhJdTX1D0h9Txm8SuOgsTv+VT
OA2yhCZLTGJIH7MjLPialOedpEs+lP8TRypTdSuyuU157ELwIJGhxr/tI3cj3+UH
uy6nSEtsg+W5y836pIs4WFUMbgmxXQH3trVv6xysIznnXxUjPG06YpMXVcuVmb9F
wnbeHeNlpnJHjy9W4lEL57JT0i7e0uXrpoHnIBSAgZqa2RUT6dYABXDni40XyZoF
tlgdGfzcqWx+HxoHYGnWYPaSP8mYuoSncTLE2P88W4eJZH/PbVc/QqroPqcgqqAd
G0kfX5dSCSLsXgfeMjDWRqxjWyo9Zs+GUQl6lcC8Dldk60IDnNWC0FJPeermjmk4
T62dnUBXafLRkcsxCMcUpG8ypZWArEI6prAHvRBtATrSfGmePb81w0ZUxRmz4X1I
+MpomQfCRnuIkMjZSAkmt2f7ToZHD/6n92emsbeRpb/IoijzegeIQMAUBmsf/T7t
D/y7EF3mDekXKGCqPV0bwhrXJxLV64UO8aE5oK1OX/twhNCDLefLLa8AiOWDUZZT
hfsWamRuQvm9BtrQWhPdcxpLP0IsRp0ru2Q5fmf2hwwvU+/PNFzGL7PjFDvnklBA
7jQn+qX6vhjYNQ++xqS8p/CiD6pYfNfqz2/QTxkxS4pOx5iKwvUwo7skjhYyhkgD
baNX0X38YQPLW5lJNtbe+YKVfho1tQb126UGh7IHmR240IfTCvmzeb+EJAJ+eyDT
fzWs3wsMyHO8/nNHtAJUwi/+Oto8DLhqjyjVSUWfgll3asZhAoZ50nfJ+QAX8nmJ
ydqJnUTrCBUiIW/CnBYD0QfxOKn3kXdHuHL3f5oLE3Lvqlv6O+m2FBHpEK6z+t6G
RZpaI6lxgFm3AqT6HD1YLT5Y/yWZRjKZHTs7asyU0XP6ZChmyEcHr6+x5I+xiWEV
+boMWbUpcBRkFkJh8X65RTWl2XqXD+W6VViiEbyzsIzWBMcVizptMIH7PKPebXHW
YKeUFbOz8uR6iwXjOqmfu7Bgg+1O+Xivnam+FX1QV+h5FU1c7NvjhJ8nmVWKn11w
bqfM21cW27nXhQ+7P+aVMa1Xvnz1jFq8UU3tSV/x1mpuv9keMMCekEqppfUilNit
jeOxE27dWFVj03Koue394MI/K2D688miidlIgNsIhWL6tQN7rTKqxytmKe60+79V
nuC+l5PTKK8Vt4kKd6rTU7qoyuJ3IIgLnwxH5lx7S3w7uXSa73/SKpSdtWP1lApf
zTJhqE3lDvyp1MoBymQ2pN/yZS2Wb+jLrtjZwNZAkLQehGmbXaJdllZlk8eVJRqd
GDH8/npVRMj3CBB7S7T0cUKnvoZNN68bESharPDmZJ02X3+9FSRbvsWwn0nYFonN
Wn98nD5GsXS+y7i62pun5D7hIa0Q2HuozezSgTw8YKcgSYikE8FCD1Bei+AzSHYO
36AiYAQttD3FIRHYYfAuIcrvd7gzDqBhWOFMAgTbmV8GEczX8G7rOrU1F2+cC62M
jCZojeC3jV3jgww/wqhAnMZGvYXVR7+lvGs3N+gn6qz3JkWEBnqi1+DIytIus/7j
83vkO+ZuMKYMVEFPtt6gc2eLjsWpbmNMTu2NeDA8PGXKqtnehYI6rlhDxgrlYp/N
i6nQLTVQsufcxlql3le8/ydXOIXYPTkpCX7BZBMv6E919nfqbmsvNu9vTgwuqpA6
HVI4Ol06u/z1IibicPjHjzpfHW8QT9ZoXhZ042HfYga9eJ6EkCYG9s+bcgDe4Ygf
ZYfCmsnjaU9/5AUboe+E/X3Qjwk5P0LWdXv7fV7anw/xFmd6klXjXDy+5wVf9i3z
5ySS0bbxddX7licriw/hXrnUD/DByGgEG/VXQ9qw4pJ61bOswGztxMXZnnpWUsQ4
1IYjPQBWQUONYpD8G4QfPy7iSOsslHrkkFlIKOPVrjq9ZnHb9wSN5giHIYFseziI
D4lQzH9eZ/Wg/qD0cLdrk0crEqfhMD4ZBA8Hx/qfAMgiifoeBuJa74ZizV7JuEIv
Ajrz7Hu2XXuQzhmIe4ly6WS5hQJkzXwI5kyP7kUKa41HK6qYtsQ9I3IKpvu9leNv
fD7Tae9jcMPSTy3+ykZLwHtLYB0t0qMcckle1GENh07oTis44K9dg/Afty7PGPwB
b/iMZdy00R2A1/lyo0WAityiK4xZFLsZELR/SmsMqHNu4ZE6CjF57kq0ujGsA96m
jYwOdEhhbXiEEd6hkCqxhO0xvwbqcRqcRKRvfec8AdXmdu/tYygLwamorvlR0ccr
qB7aQ02NzHkCqt+5X1eLcq30RD3R9YQuoT5DVnGbqspA+c3YaWsdEUvAJV9PW5do
inDeeMggxIiA5iLVLnEoet2xHTrHb/ginvQYtmo1IhPcrvoWnz6zt8eMU7IBHzT8
06kGy3ejSFnefyxBm0jla95JbwsIyBbeJpFxd/34S4rT73yUM8coayHkMcCTf3Vf
4qd2xUFSJCQJHQrqyAA8fdbNKX8DDkkS7SCKYlyrTa0Rh1YAJ7Q+GEFxund94LGz
WSwWEwesEe+7OxdeuEpWZVpqe/ONrjCyHQBW8X5rbCizDAuVt0gPyvenTsyzkqfg
bvfhddG/fJCgXVZx/5HAGLduD9E4Cv9LvutcqQZKYHwyVWomuY62K2NgxTWpWSlz
LPqqzmMfLdrD9omg0W0xolSIn9PeC+CsJQfO1zcmi60vgQBrgQ3hy3vGQnpPTj27
ESLyeNbsjKq4COaYlE3isQ/j99IpLLHLKDWbVGAGrfQ6JfjO786S8vyshHYSXamQ
2ClNM2MOYf9qzOqBOlohsHGv0Ymbx4ARiAHxeSrNqz3w2xhxgEkaQWz4jRXeR1Re
JcFO+4DdhS32lLsfhp8LpmO7UT1M/L7yvN1MrIX+1pZlUa2+Dp+bFsSBa1F+6TNX
dRuetPGLrES4CergFpKIKRcrWwD9qzFhLtpYpDtLdazxTl5cM/IFLMq5iNmraBZ2
Rkw0KlP6UATtCP1ewYJeq7451xMVYm8PNV8POPJFVM7WUkBIXzImDfiAxeANJpbB
/8+i3pJYnZxDMKGReZmobFK0UM7Xxj22up8ILZLL9DqxXMncFAY2S+cOMILbv4WR
6eIgs8hYyTIez4jSpiH960Rd/GR5TQOMtHoiDdXCmTWPNGCf6vAMgNJT1ZLjw9vh
DxvTgGGtcVE+AssR29Cmmsnf2ToL+kvb+Py5X1s9BiCxFUXqrWxscrlFTwIOoK3e
UjFP6qUswngjkohhKEzZULlhc8SqgoFjR5459PF/pHTIZkQcMheWS6QHx2DmFs92
13ufb8SKnif5juGWOvGbfG5UzXa/6XRjAKoHww6oED9MlB/xbY/5bYAYMe6tyiXZ
Hbns94TQvbD764KUwvtt1Y1GN5eJjSSfM2wZV/ysyQJn7IHVpcvVVkMZxwb8eoMd
um0u1Tq9H9TYjNkYalu4/8hBNajp3Vl32o4PFGvWP3EIxa4QzWSDXcq0IHbXavUC
5w7rTB4Es4Hj8vvX/foUaboHkT6JiuAEPZP56DahW7ZNM8Bpeh1sWRniqD3pL2Vx
nZRRjX7k4WqgZoMgm8x8I0FBWI4uei3GbiifzF9wQ7X8t1hck3WXiehhW7z0NapX
qK7oTrO2jO5wGCJcpxUlKRsvrDZcJZLplVFJtzP33z4/OA4t/2aktabL6j4s5LoT
cBjDEwtqkvhnedMsTcGAvtLjavXclWVla1ErFezxqrXjhWiBBWlQ9L7fiHbosqoz
bA23LBachyK8D+/KtOrCtRtgaEBi4PEQarYJeaZmmP0=
`pragma protect end_protected
