// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:07:04 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pboIQWFdB4Ti+DCxGQeUfmYCv9ebQ+IHsllZF3fpc2xABb+mT6aC+ghdJIKboV9d
CtuPTHKz3jdDVJZhAJTJd/p01F4ZBzmRRscucRG32zeS1jZRHcfby6yiitCOenGc
2VN8XFr9N3ZGnKAV0dvH4KFDqGeoNgzqxl4sbWV9X1g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7808)
gIaw0pPWdSuRJp6amqaUGQ56f5iUNu1kzMPBOykczDsxE3Z0mPG21Vl8dQhDjgbI
EoXdbZkaVfpGKKsSuciOmVLXNc7NHJ5fz2FrYLELyefP7SrxLlBXvHKc5UDBQxun
0VggFj+nRjupIMKbPUYPWBvNKT2lAvyfRn0R48Dkx6UxgSCQM1ZiDZTdvUalHvOo
Upyeuc/iHjA0Mxcr004C8elWe7gcE9H8evYaX9GO3fFm5QDroul0Vb54tzIOUIKI
FhLQhqAWATgjzWFZdxpvHFVxoLk052e21HoFI/d7ssmKkjxELjLs4N/S1iTm0VBY
6gvNyaPJqLjejUdEQTMNlzd9CD6dMIMW9mU8GZgw/tIxJOHASDW24FlhAUbVh1WM
tVqB0lbAjTAFn7P76i2rl/iZuuLP6HJMzilH7b3zd1Wi43juk3Q/kdu9PpqQDgp0
5gel1JB9JN8QC41GUxGk98jnCX4M6fU4yg1NCiBOhnAxm7VUrwwlxBxERJtjf2aG
+yi76HkCK0dXmC2pq7UnnPjzob56ZoQfFcPiuIV866ygEN9An3GpMfKI56adviOo
IyFB5dpZlr3vkLmEoMSRpcw0RXeUGYe3GyaWKFX35V0pPuMEzpi2IE9DI/xAnO95
Fm0mK5EbqNpSnaUpjeB0iu6m03F4OZUItf98PB56jgPgRXqJSvxEkAXrcS5kOqpI
ieLu985OlVyqgs3JpoJfDU/lGTHE0Ob0gSnS/cpm8cqV2mzrfuFbLFYcP+Kf2JqG
9MGMdWLw2fqUTOpHvh/Z2c4yZlmGjqhCZ2dMQlqoUsn24G2dsO2S9BXWCmZwLLz9
ypCdn/3SaVsYjGAELBKqJwGeadb0Fx3ac6AppXWzGRhTdod92duE8rY8N1tGP3gk
SNHpvehA0quq5TOj/WnISENHna50cYjc0jkgyD3E1xGzQuDLbmGO7eilMIvjYUww
upNltPNvdduEACRQqgjHtenq5COxYum4hhANuL+5UfzE7uPrDL2WLe6JQQ8a0quO
/kh0LI0mM8U56T8jiS8nhkbF4nqqCdn2e2jWq1YzD+oXOTiD9+zbt+vIGQI0m0Im
8aSXad0rjfWezs1fYf8s8b9CrmpvGWp6O2mEJYwwLc3/r22K7XIRC2KxIRd8bYUh
Sx6Ic75d/zGLKbIK32e0fAPw2b8WS1ZhPKmF06acSTJrTwXnrkZLapJMc+44vLTd
bg4DGUn0/Vte7byYdNlfBIYm7MAjz6VpF896BdhlPbzsqxL17gUn69kfd5ynjfaC
mFskhAwLI8Gj1BZOKncw1R3qA+M3WZKCU0rCno0e6BJiF6kv+VdF1aKRaPGpYm5b
2/PJiT+sweedWiwqaVdeJ29v+XU5asQzh1dO30ayqqdm0MmPOvSYOOBUhjND+8ua
Dcp1HArc0e2yocupckOuMoABXE7guME4spc7W5irOW+2N39yqF4zeoX/ZhzXmQSW
rEUfoXsuPR0N+ipfyZ3j8JSnElCcJGrC0cI4eFP/0mnubzMEWw/X5DCP3wMlMWZY
6w4n/izFGXpFo7aCPmk/QXkwj0mFdnv8iZaAmNVQYr44ED0ov5FMn/cLQWtmkQck
5ypwNWgloWj82liI2ytXaeqPxOVY8vnOVa10U8KJOs2T9MmFGb16hGpqwIezvHxa
Ti4UH1dsuP90L4XCIOd0onzzoDyb2fyWliue5TkKLIT+69lszth7HsIOTok/cLzV
2geatIaiSuxCX6Px2949TxU6Ps/8HguDbuTE3sH5CEnDPj1aBzryWskydNXcUWsE
mzay0ftYfOcmPmT0dhwZz+Hfo0qGwQPoDZkPxOLkqmbbVY9IaJ+O0KzDN62f8Wib
o/b3wRTdJ3V/0gnu/Uo9Cdoq7bka610Ka6t1iApQ4EfFcyX56m/Kpbq6qNDfFlqr
3vOUK7pEfW3PDZifCSUAYzyyFnHwskZ39b89ueniUB5MAdwDEnNJLcXd0h8qro3q
Lg1SJR8cFpGOXQc324gewXh/6hyFY8/gzS68AAAgugtRBfNVYfBWWyJF9L5mCC3b
d0LB+/ZNmHvkOmnNy+n76cwtQq8r/X6hOgfC3x64bJs+8WUvoIhu5cBJpSvX0eaQ
zCMWAnwtijbiIcw8XXHAAz1mLW4pfHGG3gt2AriTL2TydZgmafSp1uzEPX3tcr9A
Y+UEgHG5Fw0jheP3Jo9sC2ClMBLimcDEJVJu7svGMfD14v14p5VtSFtNOlZS1fqj
KsOjAOrOAU1hlPz477IIGnnxHhESTkuA9kZ2aiUKkp9CgBicgNlId9HZlvXboYo+
6oIb9acJ4t6GFIt56eYU3hKw2XnGVdEZ4Az5fXJiwgxhNHjFDyyPm1TJccI3RhmR
kDkQ6cHeScxRPFxzbek0PBoSIfXC/47GcgaDpYY3p2fSW7T307U1T9N7D0nKFUtH
9EYsiYcvMd6Z9llcJoSd0eHHyZWB/dfpaKHCVK0A8uVjTu8S2k37gvIAxjvaIcA4
4BNA3xocUhPbozcKzepC+BSxu9yq3Fs7Hlc8bUGkcl6b4uXtao5ETjSwT7ZLy2uD
4dyQHcCYcapfVKJpeDPZvoFy1D73INHZHy1Uk4lsEOaSPgapMSjeqm/P0c5C6Imx
hE1rTb5CUYZw7Xotl3Tmmnp0iqVFhAH1hmhoaaoa1EeiA3nnb98K4hEHo/ExKjnt
t6vUB2iQLHxFIOpwRf2XzATtfNYUN1VSKmLSjnUbLVlwhoWS3AcGTjQ1YpLfyjO0
nfvw/PAliVuiOnfqdSPBz7MyDV3gqPya3qCbD0CtiD0JCja5g7Lg9ExJTClWDSUC
XGgbAy74BMSHo8i+n6O1UaSs3wnK6AoaAXuOIhbna5na3OXFhzZgiK6Nko58QoJj
6ks3Z/b1fnCv/jYnxN0tu/SiGk1QjlfKQW46Jp2dBPMdZw0lG8I/DFXCXpCHOYlI
1GdmRjtzcMSYFKFzMqc2EqsB8PksJRcImvQ2VuDaIRo+vprvqiMtlnLYREPXCmmq
ywTHkKUkWG90ZZezxBQLRJgERLRQJeKhnB3v7SIqALySx8GrUxCSjIzW2wTKC1SR
ursKVXjdLasIRUHCo1I9pFGXeZaLTAEy24FO1kmt34/TIm0FV3UlLfpZS/MZJAIw
IdMonu5GjqJ7hKk8Uvx9n+0ZJ51czsrcHpHZuNaQL6x1CVMNBVYkF3MYRLfRRC9Z
JK6vxUVeiwn6vO8dchujSECu8DOzcJxM6caf/wZTjt2fnKIALTdvKTCjrCDEas+l
wsZIiIBihcq50z8+jM5CKEkED3WkiV65yAdTZu3kfILBi7MWTC2EYzLT7pABiT46
eAhinWrtYIwbiY8ClMuRbwkeo9GfXxeGcBBXyLALjZkCKT7I3hMZTXhovt50eeo6
LwsqsArt1JoED8yoMcENyWEYZuZRhCP2On0uLJZOM48CNQzGtzKafadmlpZH6c7Y
6Vz9unY/xJPgvxu3/xUL9GfMBCaWm+gSSg0wxfp+0XsJB72/arpy4HK9sY2urWGW
C/FZ1RlH8/tCWJk3q+y8nfVVG7R/olyDkHTGl7CuUSuOSAg5fj06vz6+qNDKAYA4
bxORXqNvKKIuMvS5yJFVraD3z2ChE3JIOkb1CVbEWTzQ+9j07KpNxYlwEu4uGQRP
gyGmKGCWnZIOKc9VDK9hRO7zSnW5+B7lnM0oaDiLqj3yfWJMulvzvdrWp8gK3gaY
Aspf/pgcmeu3va/akMaybtS8Mk0cLVLpW7HEOc8sDAlVH1kXFisihKjDtZaTQHVx
ec/HX6xiX1uTaw7/u0WkWgsqn92sCO83F02EUoAEGgVvsfGvPZcbtf2YM8cbv0yQ
g6PzbSFspMpOQW7jia379yiMjPGkJermrPQ+AKcEeD3DyljOG4BEsH+flFuNRdm0
jfRyuy1eCcVLfPer4ZtfmIPkiMZbsmlkkDugvKgXP9o6hrdD1OzzfX/wK81ZVpA0
UNCOC6sfuyhjZ6lKR39jcoLdrQhW6q1zg1sZ3tJV+r4+xsxcC86o+rIBtD4FjZcI
70WPIgFt7pUBWN8dyaPT9CKYORXK3nXx3z+FnvnpcR75EfSSsn9MmwM1B1pTGf4u
4ibyO+eiueOafl66MObgt2NFGcoiJ/e6U+N6Kan/sv+QtITTkQPwafsicghx1ez2
Sod7fOPag02NNAUSQ0XMxGYiYsZ0VVarA5A8VsmOrFARXHT0Gi2TOWjhu6q75HPP
wR+PzL9jgage5EbKZO3okiJRdM3jhmnYQgj8bLdEklrwBX320bbhdoihhoOoAbIa
OfniM167CZIQsqnLrTVZHF/6ApYAbN1wvjF8JK1ogCVtvDaHLocx3LHf3D3PDMsU
30Oa2LJpYZ115CU5Q/G8iE3KomsFWixBopFR0t1VS0VpMookcGP+w6J1ioqwMTls
tnv60rlrh1QrvA40wwDODa6tTzoNtAYqUxPRK7x4IRovxrfdQAFEPuOXKOhxHQ2P
CINfHYtkUKxv46/Fnnivj8bh9wtIS7umCdITN/LgDnp58zFAaBrbrEsqevy1I/lZ
yB1fedkDF0yS0WS/lhPtDyy1P4EwkyNVcltFoVEBOrwBpXMuVM5Ew0ICfjJS2oMm
J2SmtMdKQ9BD0DuIkoj2S6y13q8KzJc0AYfuySDq3VmStMQ9cyisopQgUo9VHQ2d
oV9/zKNiAPWCJMr+lV1Q0sZoaoIKdb2NeEpkx/+LQSa1PKtS7yTFTC8fezrVEHTj
FHYNWt/2g/Ai8cUoXxayhxZO8BPaPrb+xjGVK6ytO+quGZojTWcWMeDR60DJ5d9b
D5p3Wqnot6nlvpkEjIuZaBVPVxZ2y8Iwu7Ie4bQ4Tc/EOVoZ/v99FuaKyKdOcyb4
OIAlgej59RMteQHzZic0wvFfoa8LSDYzQY1v4bjVPVkLGhKnJWaa1Ihk2U/+Llrn
VS0Y82+/pL00bevXTQxxSE71MpbUSiRIa7yEoofbVNk62ZVbpDDezQgl7GszjFW4
6lmQyyfz3IOmtws6vNYSNndxS8kdocxf+Nx4jRq7Hw9CBchvAdjx3e3Pd/L6DOQ0
FouXZdCmRZ7hNSFIieLIreqMJFDA9jMALYzcBbwroHEUOlYv6C9vYXDoyzQzBzTs
5Y9QLZSPIuAsw6QkVDxS5HFbkgYzH1v2W6wz1mtHxZzwCyMQqFQOB4/7M2gItWK4
eEibocdZRxWev+utv7FwohMkrB8Bq7VrLDQTV4FVdgGg1nHSQs49907/7zTgPncR
2ve+iN7g1RcLt22MrXWaEyVutK/l8EXvl/kHOtg5PZzyuM6EZNTceAVdLYw/M1Pw
uMKQqBCt5qVPuaufORTzx4M0LidWnujXyU7QQ3gBbgB7qp0NbZJkkCgTxcQM2tCO
iAfwYKHpirMOQ/ZWWWNecTv/0O19I/FShXGlwfJd5GVTdP4MD6eFyI3Rfu67IM0k
If7s4I8Q49ytrBkmyWLUHMrLMtqHWU5Va2b/XeOQ8EabV7KP3eVe8ZXQA8EEodc+
AnEaVvcZOqRZzD42sNoceB7ern/wlL6Ls8w0o6+thU62PPVQDRKxgiiEBmOSQqoQ
LTG/0hUMMQgs4CoSqsDw1J/TlkYd1sNm7/h9mU33ruqsX80d9XUlRXLICzNLPgOC
gjuOlDHNkBD51rwXese1NmEbky5BmT6tSpIAhUi22zO3CmGIW4G+Bz5heFW4z8bd
xSefQ2mqZ9t+GpK+1JE2jiDvdulBx0/jKFQA0UB/h3OnlfPpOJvEdvZX4GnUB/+y
RcTgx7bOzRlk7iC/kDjOMj8qFMmrCoeSChkl9SNtJGislKrMTBeNZ0D7eWLVf7hw
YpurZhUa9H1sxdeCobgTI3uanPiuesyX0EiA5cdOHX0XLicBbrJobmnMZ+UBvYyH
Qgh/zD6dIFamw1lXNS2C7wW40HdEhB0j92T9QYmWkjAaCnJsUfOmhoqm9o+w7KI3
ilgQ2C/BT4hba+ttCnS+419KWrDfM5OGQSVlki2JfYEGrgUJl/cq0Xg9vlg8QHMi
csUAXu41r6Bi38Bdz/FjepCvBfk2UmFnZgwZdPSh+GOUPH1Nw0c6hsoCovBmMdTM
mZ9pbEFzDyVm0vFdYfd0pfbQcI3tQ/t96uAlbwm/JjXhJxQq1jf6KDcP6A+jEy/K
4UtyvAgE7wmQBznVUJCKCy/dTwDhLpP4eGt3em4XvbrVZD02hvWp1ASdqD0znyqK
hCOi1bxecnMOCxGAQuL2LNd5lt44dcValnK4/obvY9DJkUUkaoLf3F/5VKjNvt0+
wQz1AmKOm1ajAnThn4OfgytK2BObp+dlBO6nOzv8dEPo5NwKz+k2tc3FSVwAKHr3
o23y5p3wU7eZDXahD/TCKl+30Ej1wkO3elVy+/5XhOoye3J0wR4YdQoVEtunuNU5
mNRJ9JpkulHYFU60s6PQb4+eFVhwFt82cKfQ9atghW7xcwX9Zd2e05bd0Vzz4WHF
BEE8m+hHkp18ch6ud5mzJC3eG9fA3XSkD3OYsMAjA7RU281g46bcAIfWiDBNLO1o
oaMyfpEaOsmOodLEk9teYyqcycot0svQT52G5ZT9/ad7V0ZbRR1UlFQVXL3LOVJJ
ZAnanp80iiwucKHR5Wtnp5fvOOoN62AfL+XMwYuBgPVnlaS9CUvnoj81/SHUjmUp
tC4nJAFAabKkf8rfKV+abvzsIspJ3yeSBmPPnei4XYnCPIuAzHe5NAjgN1Ub6+ZK
dwhHHGeqdNh6dThDgaA58gl4gUIibnOe2YDyrV/FvQJab8puIN1Rbm8tU4U7kXAd
d/rEENDH+8d251FZmUbjspKP1VZ841A0iPL2Mhd0eR7n05/m/Yy6OBEwGwgvp6kd
d46avvnWqu/16PmeuBnMox5hMD+Up4ko3UqvM8xlxVF4VSxbF+XyLOR20xltQCrn
0RPGuN9baVmHkhgU4eDXvsbmvzghe2t3xBe+yMozCPHCl5MmE23RyrsHxr0IEaVh
kB/t4Sy8PYqWXrRWhoom4qglvMoGt21D5SxBGSI+Dgj8+ez74uMcIiSTDn1IK7cd
7mkrMsyJAC4TNnlx8SHioVzCu43L0U2oiRUprfpoEY+CaFKLxmX/bWiwZ7xD6EdT
PshDFaGnkHSCB2jOeq9GzB2oUAQTb8Xk8pTF59kCBThT1P6nQnafA8cxFcCBU/N8
Wgp1CZkU0tf4bR6FqqAJJrDa9AsJ745n2igYkJfxRGUJBYwynklaII6Mg9lwGGcc
+8nyPST42mn2wuL+20FEW2tXBffw6aOiDaO5Gl3j82VPdRS4CjdHP4tbW2VvTN4D
GTOzurf85hK05YFMvjoRYl1Dq1V4RMbeHMqbbY9nDifItz3NOEnkDXIoRV/BUqkt
Zkk6kFpZeUfk+YmgpnduYpBMuDMZZOKq84YV/FpG/YXyRhOdfzpSCAPZqO+ElaZ4
v/HGriObIoa+4H6KRdUxsJKllHH9w/TmsIqZN+3zdOCZ4CrjTs04sG1gzeUoiGjH
ZnwnkpD6cDcVR34pRl3Rmh9i7Zf2tMJlo3WmeS5XqcuYZlq0xeVKKyGAP9oRxXAP
eNIqt+741vHtxuyDuP3rExqUN4cr4WPNufOyKyVC2R9Pw61nAxLXpp0oNi9si0op
GwGoTySnl3UzRsWt0Vw64N/FB2pgQcmzU2h8BpopgZs0BZ3AKUJUOPCURiJ762fk
KulXZa9qyZ5Fv0vQjZhQeQOlfal88OATLzQ8FhuhT1P+YRjjm9UiMvCwr144AOko
uxOsZE8bhoLyp+2pBSOGLh+MzLAP7OIWKeFqGWKsDYhOP5Go/OTSs5ThRw8sPBdl
3FgyW1NjPMMdHQxGlWFhHB4rYWl732qkAuLE0bOX1R4UwaX1/S2Qf5XBiFrkBCW2
fM+SRni5Pn5tjRA+ORwJZOdF9CKvBYvXF1I89/K54Tm6hrFIjZOOqMG+mp7DjxBj
0T7draMyWAX86nC0kajBqq3t0r5Ri0mSGrH3XJLOeHzIE+HN1B7LsCSoq/6d6pym
uAfo7R6BIFEqCApVEE/M1EKZyY86fMrl/xvECDw/l0b8Nf6ZBQrmFn8PxNw3wtpB
QOpiyiMsEPZxqGFJ6qE1Ti8HVkVsMBcPNkP8SyL5x8IX3mPVQH58Bw3iWEPRcyYd
d3BzBgVN8cMcRsvLjtqTF+tduYM/4BqS/Ztz5dnGhYmnluMsfDXz/F/uHOQR15z5
vVt5pj1oMpHiFbw5Bd2Hw8UipztY/7RRBCwj8QlTG3JMLA1oGeBW3uvPEH7mfOgT
isde2tcesRadlTyu2NS/PvWvH0Krg0X6fPcbq6TWMbVFDWb/MyX9KciEoeTe2UfM
4ED/oXAE1OgRXR+LOpjefMq8mmmJlVJ8ZnKtm+96bLw/S7A2oqI3XU6LL0uJCMab
h7WhWTkKROlJdvSJCmjiyEc/uU4XhjPPicnKrRZ86dyPY86TslLNIVIreAS04Zf1
Gf9wM63nnHo5Rk1ie4FzpC1oy4/YFhIWxFGjJhwqALr5VZvJ+i/f3soGHwU72upW
+Ah7E1C/Z3ryuNvWcZXLqXjGigaCgHobENolpcEZC4j7G9le1HisuBnzKBk43z8/
40gdljeVouoZcY+RPgIE4VJJPYeJT7siUPhBNDbIJzzbrxnkERrcHISNZgt2QUPl
7XS0EhfDPSzRrhpiJX5jBtfLOHft74PlQ0wkWj42sCSYtzANVBheGTRdFLxymAJt
5kb8VkgppUrX8+ZXfYIiO2vptVXCiQ3uavdbsRT8zTRBvBJ2K0Q5bPbbY7hzKjxf
tQERIUJTA2HBw2YtB1ngQjqpp93dzqsnAvSOXI78WZqD5+3W/JG/3o4mpiqCDW7Z
8PaAN3WSZMTaJpX20HICaOoO8mZCPlEUbiHaLHX7LqgXG+i4gXTp3pPfkabFO960
wYNiXrbwgb5suh1u3v8fGI6/HmUif7gtJE7jBkC4epJN/2/MKwNvWkKWMlWQDGC8
TKl08ANjYoqROyq+vRQX+C1Ukacs13EK05c0ddHrgQK7mjP3t6Id8A2xSkI1gpt0
UoskPF26mi1o90ktAjTOs+hQT21XNmdfBsFUi3C0xRaS6BU9g63Sq2h5sym16eOc
+p+5KQJJA85J/umxk9cUc7e6lgXCWCJhhEkTW0JM8jB+Wq57dF60r9zsOY5l/ymc
Rg/VfjnIHvfhb6o8FGLMCa5dfOY7ruJ6gRgpsOHa3ZT/4003uUo+/TXrTbzoHa5M
G6SGizi1xKwE3Zt75f80qkQr2UimSO9OZ/+wE6ykjQUPZpO1WCcd2JAcn5vJ2pE/
zUQh8ydtm3HcBbKX2C+6kkCbooqnMfWLLt3gXFsqxXCfGVGNqpikVUMgw/HhlttN
4JJwTm2lsodqxke+8nxmcusJs3cSzRj8KrSMiN1m3uMY/UIFVuksXCHVNdki/Ye/
0Ik8xY3oOtnvSld36yMaYPmmaBVh/lVjgV8PvVj0ELKrvFNdsWgTAUWQAMbHmtqB
klihXgPGZ15SeUwLN7U6KtcWqlTrU3ylzZJmSryPebAsW8bX6/0CaRiwA/4w/xKq
j97DOGgd7LVquqo+G6tE22/o6n3GKpg6JgiugN73vAGJoLqNkMkmztKy0TnNjFrx
v+jFXcJc5pqDrf31SQ1q83qxx642bMR0O8HYhxcFaqBm3p5n8kBhELX4hH9SYYtg
tV4JYT5Od30yK1fXDXnfIv8i2XR/oR7mskkd+HLGY96Uph7y6byEhweXtgxjG2nJ
dZb/KaXGUiOOZiUpMRt0b+K/v3X9iKdPGZui+ydJAWR6ZoWMjWsrShHpNSMH1Eul
vWOB7kZylfVEI4CrnCfHDSOj75AwbWSa9e7E6sg1GjZB2WAGjERIIbRZUAyu/3La
xckfbUvvcvvIOGTVMtaD95JkPTtrvV4gN+YnAO9peuD3l/WqAYnvTLr+PaBEbbVd
yBgge+9fBRUgGHw/uG8w+TbRg9bd3na7J8yelug4996uM4lsPTRpFVNfGpygEg1/
ge6vq7+ci4FTMfG4y2OGEtT7sanSfQ3+NVCWpAaiTeiInuRixJ+MARo/gOIMz7xx
6Nc48XFs2kAN+gGFNh7IiJEDTpOxUBl372WG1yX1qXGxxMdLD4Wzyu/0MZN4mH0q
jetqDkPug4QUpXu6EZvLViAGlCc7g7/H3nq6BxJVlMPD1HqzgtwVpVkUF8gCYPLM
AlT2q9rggt2hj4OkBKFl+b8k09f3ERPnq7tsgQfA9ON4DM/b1QQ4chwcVjjeqbvg
jqJrLp8/S6EyFSZB0R9HQpCBsUgTLulYmaQ2HqUYlcxtXdbXAaMA6i1KSrcO2D4U
cr77+ow3P15yRWxKC4bQOkHIQLt3qjhOcVo4A6c7wFHceBCT2+P73Q/7yggqU1dW
+lpKOFW3ZOIT0tAyMQJZ59ONeKE3e/mnXnsrWwJmeK0=
`pragma protect end_protected
