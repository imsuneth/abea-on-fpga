// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:50 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mdY8YVLax1RYn+7USodbDSjdNQwNw+70jgdykG52YsiqNK0JY7hhkEcKVBFxQq8t
roLFTv8WzXy2H8Q47+FR0GuYs6HmiS86VsvF3W2PstqznLFN+47NwJySzrBhhvVi
VkxvMQ3OdAmyxEzv125LZbWj/LlKo+PHhFLNVEioXjs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11536)
vprq11b5SiV+0i3PKYieJZ6/Mti4MiUqFjqREHjf9iWHH8mSLYuOefwdo5HT2G9Q
Qe/ULAeGJoYkqfUcjQMb3JjQUps63Mx+KzBTkWj/1oO4alzxZeG+wfeX9BgMJsyy
oEzeJQQJgk+5eKpkNXGmQUwg7Drqf0FwnLT17la8cK/dyv0QPWlOdoVE6SiBsB7f
Rsk+wfhT+9Kn/QGpdHO14znLaVLAT7ZioZV8S7ZDxJdybkh60GlvkxxXb+XpoaqG
k/84VIwInFOYttwL1OXTj9wQdHLLDDnm3gt0jmIa7ezB6I7cEgIgYmprwtC8MfIN
taU1oeHuli0sY0huHoN3MEzwiyvYcF9oFBai6GHbTRYtUPdjdsNjewUUaq2wFaPB
jJb8w+NJCDjMzgSZNREdhhp6DJnKY4Tu5eUr6cMFxQOcccpKkUaHO7u5EBqQx2O6
krL10eg0qpY5cojuTF//4Umi8Dgf6tht+tAPfP36jTkJY5twtwvQtRnruFMfUSB+
d3t0Wt+qUXerScJIKRbbMyO4+BY14rUucBVQVKDCmT+a7WtbAmsHH27hqxPlmeyK
pUpyI4WBwSHb1TWUOdiAsHAFVFWryQf9RY4k693HQSlx91EpfRhg4yCjoIOUOnbj
50gznnwkF+jvhuTFUuk3WfKIIxK80QtQPTXYN0/cIYWEVXwEOzt2VOaE/v6+gLzC
66l/+T8y0FVrKfNTQSVkhqVAgwlwyslC2XoiZdZQMh+N/sbWzWRtviRxx9f8I5t6
hY2RlgStTbDZdo34QQLP7joZQZCpQJL4t38V5UbCvDJA1BUNATEYtINxa26aSTKT
PRUHGL+KHu5MdrVLeBDn8qcb0YjYWV1+d3RGdXPkiQv2jk4pk6SaLAsDC12RW0SN
MOBO74c+jck/JJuAYVXLkmRgw18m/nb/URcYLWHTc5dN7pQV+buvEvak/3yRUyIn
hQFXtp//nUS7xk7i+t0Vnwr7cUsHsGtc02K4cPPS7RjR1uBieN5J//RsBWQWLeJn
OEXJ3uOUZ8wL7Ba3PcUxWVLjd6Inj2E2JscD7Vjes0ZbZhMtOELXnZAZnm3e8yEs
AZR1/qKN+Mty/wpb93SB1msePq843rggiSgI9Kq8YqGycHXqgDgoB5DSZMvX1Ee9
GqTiIhaP56hIa2wpndLjF6BzVOWjYqzbmUcu/NNtPYAF+K9dCSUatXi5nwMRwD8d
/FWjiVv82LUM6hin0X/0JQ2lhZR1iZT8ltUGig/SXs9urgatPhGecSXglMzvMVZ8
kAlQljtpQ/lCOiD7hQUW08Fid2hP4N0HahThJP6i0g/1f97/7A1XFRY/t71/w3ax
aOCpFQLMMrQ8pK1LsGD+gi1nWSc8OBd++upmuyCaqiVoPbxzeyQKp7BjNDP7mRzh
SPAVUQEnECMlSbKpfrHT5Gz68M0dqtb2Z1H4lMsQbYGboMtXvnGdLDh4hpXDF/ZW
m7+oE7HBL+PHAVCOaVYoyf+xV4A2M+HDX+RjztJnDGJOasAYd1/6ScFIvg65zgFV
BQpAnFTuFbjwhAJQGgt+fig0wrpLo3Y5C3fJ19WW/3zk1NsT+FmKv+mj1VN0Cfbw
kher4TNfW6PlafYP1fGKaqoCfFSKGNV71jet+IvXLjzDKUhuRsKhma9MK+hk0Uhv
evMGQXtfK/9wjlrcO7ydtaYTwvqs8Dvstem7+aUjrK0izEZ7o7zYxM5tk6CmD0Vn
heH4YOXQUlCsxgIjQxOs17F02V+XLQmVJLyA+Vw34PZ/2duOpUp7K75yRIEPZ3b4
YMath0CM445VlEziSZsjrIZtjDzNs365ZAdpHOq7RqVJcw/OV0m4Bbe4I69IVWnz
ePG46nu4nyBHU5V7Vb8Oihsh8Nky9fANc/gSBdP1zb4TMqtA5Z4Ey3VknQcTKICm
h7ouQKSCo/11noViFPClnGW4SjH8Aqn7jfSPlabl0GDohEVVPtvDTtMwa8axPm1W
+IkE1WYfwEeExFy5HlaHqQgUlosMtjlnVVElCAoaEznooe65OvL6r5nMA2CEsw3z
9A2oa11rJ0XFb4Kw1KBuzeStyo89f9M856iQ6+0GzNiX6auuSllK1RNK0VapZEwc
DGTegQPpGbi9uo794XGMzV7lkXHtx3XUFX6Ro1Yt3wI3TayfW/IinsACSgVlo2Bt
mIGxuw/sSftqgO+esIc2LxWnoGdn6G9FSk2CGMt/UGX8WKUAdPcxF01iyyWMubXr
azrvFD/6yjhvkcJhb5NPn+kedILllR15C1L6VKJmtefnDLxg3sEsKALN2s7McVrN
JUh4EQJ52kDHtlSGrMXB5lWjWqdho0CL7VdaQtkuvfHZPC78LSlRwuWqFQCSNKxB
7fAckbAaasj09VG/w+WK1sMTYGoFBgUghiZlgYiZhNG1t3J06+UKngFU/NoZ2NGU
bWaGYep0mGEOH9d1/ikRyAsYDa6GbRXdnvSUWnrFFciG6A5u7RZAL6yBzhrwDSko
sxaLVXmf2B2y+v63B1sCmYDPfnhJ1Z4ShopnoGpuRsQcHLiKR/waHIH5/JZGhT7A
RMm/zJ38bi/6PgJsqFadvJFlwUW/rWnBB2x27pzxGRxRNhnIdXa14Jyo+hOWXBMu
LSpxSpn82tij03jMt7OdFRr6dUUX0GC4mCrgr6bH+CGrJ6djshyhPsDKqUWREHsh
mIJF0lW/qYvzFrn+zUhwdX4gPY+I//094E1vtx3vnQwH+zBZsNBTen+FLINujZG4
Q1Xs+z3GVO98xCQZyStPT7CpjH55lQNs+hf5lwm6mEY9uQFfpyvcNU50PayBLRSo
96OCCPVA4UUZ/F2HuGoq0oPJZgR5sg5vdTy6XyyVwytcQwmGadDH0bPAbv1nXnHG
NPoVvPHJoOwi4rjuEoQvL6gyWvkAjbagxmklK5vRlraic1//5q2EeBuBMu2HljO+
Rc4SKVotdKEbUC+cVEKYCq6UJsiTHFEDp9KT1SbaF2k6U3pe6Wuc7uYrxlu+7yQP
XAqhzkQm1D0/0euTCRUH09kAJY7ihJ3vwGG1wyhI3XTCckRVoyMwNziWnic0JlSY
xMJDIywysIDqKgc0q+BA4Mkg+O1BpiszRT1dKipmXAHgacfN9VvYqnNlflKn7frH
oA1bhOg9SDn3hJUeQTmJFyLPh7MOQbXL2jh7OdzdXUABHkx2Fo/3FfyEz+5CkVLW
LMlo+XLkgdT0gBQQF7YvSoU9MiwWte1QZa/pUF0q0yRS2myzuohorQKvNZST844w
jnm4djNks+rcRgpDNtkb5dNnm6t4o2D55Gj4yMZPBVL8YIQgV5gKFP6hgnkNAsT9
kB2upHrmreiOjxeNkAi070Nd/30uARty1Q3aTTQGt/O8i1gEH4HHF/LGUuEQUxdD
8Q0j+4o/JB4NjCFBLe0ofxCac3VhMxPDOvq0pUBoephkT52WxwFwY82JkEmWCEsF
A1YiCQCpkz1uylUgc9tdWzFnbtUYCfLZJhvWyEypuNMnOAYFlvq/QvrGdHvf0td9
UwwHV/N52A0eS8UK/Umogm8MXMZEg7g7Y18URcck0hO+L1qcYcitknFJJfP/s/C6
yUlFpuMpflI8HluiKEVXTlY5iBqz5GsHFpIjgAZ8gK14pCC4Ss6BxDnqoBZHXugJ
zL6jll39/XVTbkMu8APuFySSOhMPtWcdongx00bQXf4GUqXL72x4Gm61I+j+Oaqu
SX8NSMBPijDeEgDrlHlErcSn++Kq9xrIKDuYbSTXIa25+azFgg9Whk3ZFM/pL+c3
/ehT0flv/nG5p3AITnFwAhtkn34/ZfVx+1ojaPpLPyOnmnZzpLQku1j0zhPvtdbp
Qk1HpCGcXiCbpMlkVMIaDNXb7viUdMdSJ1sxoAvXq9+7XkHb//NdaDXPhrcH8m0i
Adm7YrfW7HuZ5eOUvaj3lPAueVYDwuYCsE6X5Jy1deRq60PJtbkj31NrKXFBYPE0
SYXC+tSA0r7HY9eZI+wE1fe+WlHL0dG5b/OctxdbyFU+zHDmGILQWl5q5cs+YeMZ
zCVf7OvkVA2mskbZnktIWP+5ks6EOTNmqHX1kzGO7+vSItSmWD5ggwo4vSQyZ0Yd
DVR5VxnvT0tMsBtnc6yEHGb7Q5HmFIiwVyw63tpKFW3bpjmx0JfC8WWkugxVn6th
W62WDl8M2mQoXZ5MRtFgdCEOBdQr6FZcoljMSGb4RvBDfZtAY8ksbzPI/JF33zqa
w0nwwAnQXqycw6Z/DUpnTr/7nRcGqhEqYjDs++NN/nI3X5pCWqSsDBKkEJLaSR/L
KxfUz27/m5x8pPsfTc/nJYeng0ObrdrIDpV5ewcX3guVDMscioYQdI/XEDk9F4ub
OWsL8SBJhKzAeY401WPu5aVbiZ+G4LVWnpdAgh0GvCA14ZAzunb2rxoKWoF+y8az
AbKa5VzAPoGFsajCIlHNEPO9xqLue1s2OChuhLsWcRT745NADIFGrV59ZK3ueWro
NxdLzbzR4qE3EXsMCYeK1sL6OlGfvRAhevKu8FOqZmmzuJi/e1bTxO9PzP6P5WfO
42phWLUQqRtmPsZEElZoGet9OQvoek6mbCbWas4gi1v500i3Uuzx4p//PhxObcI0
UPtM4xijrOT9C+6/am6hN97BfRqT3sr4EKJ2HgJgmaOjv00h1SfG7cFEmGtKp6C5
tCoGkcaqFKjNPbFfhwqhiSw6NWFgLa3kb0FIs8zNLvpZno0oGk+jGV4fOTpLwrrp
6c2H6dngUX75+3a9gYZaLDD1JekXWsNAc33bdMyhQ9AETmbZ7s92Gf+3wGATM0Sp
hk25xM/EqfW3bkWk5YVax5ta+jrdH15REf0rilLnuo1s+3riWBLARBIZYRJvBPhy
UR7PEbDon1Y0pIVIKVoEUn9v0u06Vh32+TMsv1zjh2VLV6+O1owKFFvbaqxq3On6
yYKusr0QXA660MbCkK+oeaNKp1KsR5AdtQe/w8eyj8UnYu+6A/Vy/spCyunC9kRW
4rWksTA7YqNQU+7pqRvAirVdgi3V5Y+TH4HrNobjPvOOVAxmmwAmRVpC3GGl1ZPB
+yFMyOPWcssEV2tQKfppQtRzVHyII4g5TahDYghwYxxvilwVQtgihxnvgH+Xdscc
okGjOQY8fkORYiLBI6RgC6O1DsIz403llIxcu5gxa5BM/yEH29ghk/sl71E4C9SC
/pmr4jMeX/tZhszNtyGMZ/EftZYwg3LI4YBzF/csDD1t4Gzvy9EeRaoV1IF+5nvW
p9uMSWG9B8T5jU6USXkbe6pc24SFqFKjnCLONmcMF/bQnjBjRPhkKNAeNGKy9Dvl
xVfRdfZlRtnrVbIJ6k8t2fl7+zmD7KoxGPkRfqACjRHwBgd5V1vh+wI0JTj+4Mt2
wb/olsAlv5THQeySJXoblVmJ7Tpp5o+0e0AKPkQo/AUNLtwED7u7gkrHl4pazuXy
LajEkNtAmV9Q58LlgJ44D1PEkGH3n2N11TO7Lr2+vs7rNgQTniVV7NJymh9BkOLV
AL53aRFIvhxaZAppwawFWpzQhYBxyZpUCAstVV3DTKSav3Z9Ig2v86ytEL2AYUzO
R9E8w2G1P0OTpiP7N7SHZgx3H0YNK6UwSui6VxE1Ar3IaWNGJLPdIx5OOvcHo023
30OpdZWf4UfF/8ACTXe30VYe3OI0BqwWPtjI4TqSTrAJDz7m3rNh/QD11rbwNXfw
usV/ftnLWqskbdsYO2I1d7js1S5yFgIgfePDQzsv8WOXh9LyfVMB8mTEH6NHAP7x
Ace+a9KbgB2U7C/32SFizQexJTWpS5dUKN73vQcDWZZHpBrsV/sE4Mu2ywp6C/9s
WU4K9nCmLGmQ7QWS71WvYwfUrruHNJRrfwZ2iNCL22HNvVXD6uN4jhFlmFhAjShv
zlpGwkAVp3ZDP8hDgG0g6eY3jmH+DQwAkbJj8widjCvxsXX6iZVTAhLRlJS3GQyK
6Z3Q9u21C+OaetOgHc+hfa3pJ7/8A3ayZS/j2g3bziDrkmZGnMl4ZMAlpZl0lPwZ
fi4ZRsMMAZsjm16JeaI5D6qeGMLVyJtS1QRLo9f6YfEPHGD0X5Njiali6KTjtG4S
AP/oXp72LLF7uJ8oCrHsaOQqTYoG9RpejH/6fvLAv5s1fFJzaCv/upgstWHFc2Qo
8WjaJdcOBk5lMfCKVCFdfa2we4f8UmIsmxWaS4gNYzEq870ww477G/y/TwdYOJUR
du8w/Df1xLNG99HqWdHfiBx7f9wsXWZyTjU13zhvFVC31FDcnSwp3QiG5fO8USdH
sKDnA89Mmw7B8dVPNH4uFxY3twMlcjBvg4dHB/e7Xk2SVVQWg3jpDQqeHSK7XMN1
LZvIoSwYuL/9yz0Cm/9GXD9xwnB0hIN/+CS5KFAuD9k4oBjvQsAibrcO+QsfOaJ4
323qtOpgGFysWgi7r/8LtnEbOtKwiy6eA+/GSDs4HbcdeCdbb4+7R6b1H4PHEAGd
R6lwWP5rJcCjX9h2bHub1/D7MQ6T58md5tyaHdYVY7XazfyDl4vuvyi3A6Kdl7u3
7yDaRwnd9ZKKVe0Z9u7y5fJZgv30F5jLUCgVAr8mOKX/K34VoJuKkmRqDvmheOM2
isOna8zaHXM3erw81B8gIWL00VyreVTg7TN5mOtf4S4Q2HuX+zTRvx6mzueqxz4u
y93PtqM89+RtCgh3ebAir8izWEnU49++ERQXUAcxMdaCDPIrtaXV0tehOjgTS7b5
dN2y9fjg75RUAT1zvxhJDGU3XO+g2RHzrvV2J659/0rlmBRAW4Mfxzc20xpecPsK
f7mTU+rxUS8ZoVxtOnsv+vBvLsvsZeoFP4VziftVHec2vIcCVn8JHttONLjL8VD2
sQJQ+FYInqZwIjjT3IlDeLXQxn/CSXK5GmJtQXsO9Moq8FkMWpzrHj2mSckO9WQh
eX/qb8uuHMJFY8UvpjjqJcn5TA1Aa4+Xdq2NNVF9ll6I2mf9H6fVc6Y35xumukWW
N9VG7oGopWc4sU/aV1bLTYjEERBymubghVuoWrpfSfTNcO0GEzIkKWT1rj1x3DQh
K7D7Qqedht35BmslmMFMWAaDQT39bm5z8Ov3Ls35k7bo3i/OawbdRFIFLMbmvad4
i4Y0ImZQI/XS/QyFYu2yDyyLNY0JIdts4ftDoTMlRSpJ0IuMPy1oLwdVm+W1QYPj
/fYJNJ/UemJbUaottHovsEJA0fy26fXsF5K30XdHPSovsa9dtwYsVXXaui10aKUL
K7CxeHGlVN/3Xva/H3eVAfFSD/nKjEu+kuO9/oGztC1lLFdD8l4WD30QCAtQOcGW
F5WeHpqh/lA2FLUIcRPH0YXmM33FoNPpKXrUh81YlI9XclwRAFqn/Q27GHgbvCEO
yjylrwgsWqGXfE6PNinc2G9YOrI8S9rtcvEiGES8MuQ2o2xa714SUcjlZPh5O3Ll
zr6Tti3RZNvD4N9iB5szqzJXgqU2XSjW9k0ubyLbhUvWZIHSHh6FkcdyAlZjaKG4
zCWzYKxfqdhzOft9p4kBqjDAJ16GOWD1MsI8KFxVTLoHf123eAY5KdN7qiebAaDr
vNMNj+qwvT2jfHTxmVQCjgh8nRolK2csQnwu3fDVDE46c0trF8Ht0a5wcHRjDjBM
qDNvylwStWUpKS7jj0NRy73an2mM40IqtxlqfzbOgBdhmqStEhfXSsgXzSvpMJF5
7Tb4gXD+FDF75KLn7qmTCwodJE/TEgCsVpR36QUAe0YwKHYCzrsWa4H1whCWBvSc
cbamepzndv2lx+itCBzyt65sR9yTpaY/MIqj4clDvt9BlMcuBNtRyMNWOHYe+qlg
4DV25Sg3Ln/udiFAVwpB8NYDCB/VU+PZ6ncczYlivT98tHvrOPwipvaEShbtgeIS
i6aMWqg5SPbi0bIQn89hHHWRxbKSJxrbeca8hMhHu/x31R3YI3P6g45G68myQX5B
nD3HvDHRgdJgEkEZr5+d/piUXIIM7RBieMOH/9vAVzvv3M2kBMQA2gqc2L8h0PNQ
C5j5fdF3UQYbHKDnnkBpM62z7AvYdlpyhZRr3EBar+yEPe9OexwtrLXldO+rUUOp
hZLpjmCpoOOFEImXk9zz7dOBVNBQ0dN9+FGaOOqxVxpKN26gPQKglPP60O2j3ZM8
4ZDgrpDdNrEKEWCWB6QWxDtLhzxkA4swwHp7UKaFDuP+uBQEmi+v0eB6YUekY2JR
FRkeVMxWZDhr4DPgg2LMKGoyeZndXrIjtXpODfDKlEBtjb4P9cPvNol3gFRti4xe
mktv8Uvcb/kNElM6Emc4XHcomzl7bQUvsF+xz0wzs7efHXRm9lbKwB2TCtmMoG4o
VTJw43tHOjzX6FvYdSzNF7BK/XV49ERN9G1kV7+0okkGzFQPgcTek4C70BJej/tF
Dd29XDM/WBulqrpJgGRU10aIOYwcfwFX0oKFusdDYVxzfEnt8i4LjjiRkfWBR4ot
KRnd77HCtudLyOr2uK0e82ZCG4dlXuss7tnk9PiFmUsk11vwzbwp5tP6HQrb9Vyr
ADMGDs+Bpw79M6o7DZkie3kvcRNU/FVPP6v3GK85L7Gj6GuSlWemCi2oumfHaHff
N6ycq0PogLAlXr3O0M4sINDg4qDxpHsw8aTzEQaOfTUgCgfTSFqp9qCfAKy5lq+O
NjXhvsTUSYwPsRnv7ib7+qCPkMeSbXkfdoy7bPWkzyAJWbYMByuFp6OUIIFZhegO
sla9Sl473XbBcgb4R49Td5PXB646Cp0v4/r6eTcMOwHLrfm+qtj302v5kW2ayAgN
H3uou+xbNs41YKOV1PMeoqecc+uUDVen+OwYDJ6Qbsj2fLrg5v/SA/9CUPBPfjLG
fNZUB8jNgSb9QoVuOSEm0r9qMGh6L3tFKtyt+Xdqr5aYxZKKX0D1L3eu9PicwiO4
0DJuWtzlgw/degBlQZ2qmigmSRSVtFAXcth8wuuotNYwuJynLXvTuZamBnLy7mZ3
tUfUSWvSeGTniTvDyDZ7JnHy7gpEKc8+MRalI0aVivDHa0Dh58u/m3bLox09Oy9B
kjWdgoEoxvkjly+OWkR0rFNJGtHdSLKLM8a87YmhgEKTkJh34brEcGIEhI5DyR4D
0VP3aIX2qoBWl8YavdP0ZW1FjavSKwxiVgsfVIJAWrMfZD993S0YoxYc7c2iEGMn
MNJ/PTg1p1jGLXICJK0/ymmpntZLYcl53iAaSwU6h6pHQBZv1vxUzwJUCAH5sXo8
0/7M6TIsxnEZ9BGzoSFetyYnOwUp6HWEAicP2VxK30xPeQ87soVrmdbUnUE5tMLb
hmtD6dmvPZSBH/dhmqqUhkW0aoGV+Uk7Y847eFzQfaNEUyCk1JTaR86wvQtopRu6
mRbfYCY/jBJCQHjtLsWH03h9lDTGPz8Aaz0tfJIhooBDSpgVZxrL4vOaHQUiQqa1
Tm9UFD2N4ARnfRZVPESSRZ50ZC3vD+IcmvfjTgze4ylBKbAhWOFnZFZRX4nRsIV4
7gyHovXo8kev/lh3reN7Nf69f0AArwUbxwSpGuZjRiv8+qPnYpKVtxG/zTMSdYB5
/k3DquFP6K9ntjyeGzYJk2eSFkBTzMzDPfu33hQumo0csCxC4JtSQOZrxSpQmaY1
IRtbUoypXBqCBoBxVsxUtMUwD9zmfMjopuoObfCsoRLol0omCmGFbBYh8a8HjGE0
Ki96+DzM9Hh0/3G7qkFbKFNLHTk2nBcI+5KPEOah9Ye9aXrTiX39cyLDjD4rXZIz
TBMyPeDYOzHiy7QFMsrxtyYvzU7kq8m2/J4vrvvLxbIVVdSR0J9bHuWOuBx0Qox5
R+7s3C/WAD95XyJjW6uyYTriYWF3haa45FPGrb5JvaOoiL7PNqOr6ns9AETjSxwk
k33MNHcsUEIEJX6HlMcUkDztz+y+yih7mlE9ouHaR9KMnNdUkyPzYQ2ECsgLzDYf
4pz4XxyEx6+O0gkL8KwfGZ/lXsK1rKEInhgHJwxfBZN8kCc5PmKCp3B81cEjG6KY
CwXTbJfq31xIs1MJu1hAjd5QTyRt2QVB0y3XUTFmqpukWUigxQV4lIk6dfsTKlqO
/VwyT3Xf8PH8Zi9wKF/n2tjnEpIgUz16S9XGOoDg4GEmQjw0n6Eyy2498/DPibyd
5TVLfdj//jQ1fJe/WXj+9lWgtkloyE43pxyJGDwgYwUnHW0vjml65wl3iz9FEGIP
DObrq1SajSjTx4Aatisst5AhfkjUq77dc/LTgODKVy+lg3qD866mlUudi7uhvebn
12kvUTdrB7/OQiiMjh43h7ZE3sNivyxjBDV5B0CNt11kSDAAG5RNAjSVZVAR40x1
+xl9aEI+nhmFVrLbNThvmnDc0VUz4Xv42+2vmAAMlyiYuF7X5mAQnDNeY/5NH5I8
yKOWzsXTcvFe4DFVm6geOVVXS0BdAcdCN23wzXHwG8K2QIYrd1ytq1tisMNW+b3H
6Zxmm58DIKA96v6/gKNAOyezQnDGvAkWv+LBmSqtCeML0wYZOo1/qhjl7jFl53i9
asakUeHeC6F2ZZiPB6Ai1CwIRT2Ex8+2+BHd4vOhxUn/4ANJidlRN4IgZbM45yRn
ZKVdogmk1ElJfba1xIiNXPB06RZmkPppUzPvORizv3HtJYqGok9uZqqbRXs87CAp
TzHepOM+dXST2yF5bX6OQ2zq96+1MLonfpn09yLrLcx4Z0ZRSsK3sn/1gKFAQPMJ
wCQJKyNDq40pBmlsoU4/OFesgX+AH2mMYMSWtthFrBMHiomz8rCsv1qSGfJM3QGw
sbN218Q0U5/LwtQnrhOgK7CQq5IQuqwNOAK0E7n7XTv0vefXnUZ3UmUFVmDEfBQ6
El2edfq/6XVzkQz1SToWQOOsGbJs7qbKs9r9quBoui8BDHvwajpuJKHij7H9YCyG
6YmLjXAgElA7zIidqnzgQyWCoiseEjXesaT72A0t74Vr5jxuCfqWmp/9EYQWeyV/
PZpC2k43+itnMcB7CAkUPgz6QuW5LmOiMVI1bgWds1gIbO+XuidiS99TNLgyN/Qt
Ih/pnivnoGAkmWa7Fpp47OzyTL7hDuEDUoEwdVcHJN9z1RPv52iadfknU+4TB4a/
NDH3VKUxcUjWXwir19QYx3mo4BUqDx4GcxTAY3jl7AxdXMftqqgNyvJ3SAJaegb2
pq5XgPiPSCouFqPx2eGbJXOsp9bGmvdZH8R9G4qkBO4ElFX1ziT1p/z4lOJNI1MC
8o8xObGoa9h1o8x2V0tPsyu7K/yp83RpKuyctSwd+QK9aVrcrO8SkHq4yZ/EbyDh
F051aJHBsD17Jvh0u0FXjG5TYIgd1gSsLvuarbd4Tw2Bg9uU+rSM3EVo8xfhalzU
8zr6rMyxela6YYyBPYL701LFyVHeybto+sFH0safTFtNTS6j9NpNdNPmB/aYTqFA
nt3vfffjPJ23Tbmz6mFMAseBvs+ij3V8tQQCk/6YEq0nMypMUdPuTQT3DlDW+L+Y
jBYFuGxi2zvGQNUnda7KJbxy98szz4wQEvbcng+Us800ADSNZuQOefY+M4ock2mZ
hyiiUqFRx8dIeL/frRSP1L4eM/FuxoVDRbmpVA3ujAtDHnF1u+jlByjOeegGAX5x
5HO+7jp4rbbbN0KC5La71aeY9dyBFduQ44TbJloG85nCLaVIU1e0yOJL8K/0FhJg
BvUfCRl3xuz/BMPlArrmxZiS7buroXG8ba7NNfMYgd/4rYG0PK+3TwHPzAhI9JOm
WR1JLGC3wruPh8zBAH616pDJp/dr4Jyv5Tq+l5kpZc4fzLOtJ4VdLM61r+ZqdCEt
raPfreQqFBkvdlGVSKfZLz0W/BChXTxJhsq5uIhkB0RM9Qi/hO4JjdzjEQUjXQuj
EIjzJlOfd3hB0sFx08TBxlZf2ORda6vg6KQQr6N+bHR1qTy0zW1HTf9Scw9d+x9q
An4/Jvxl+reQyQgCYd4Vdocv3CHwbJ/X+PR1Pc0fdeIy/fYt2QFws/afqSLNoe6x
/o0M8ICtCq8tTdjMa8hqXRJ+YdFYs0sO1f2drdIK7Pe5wkp5tWGvss/JBSAbj9zK
yuvEnOhHKjOYXhlc0BHc6KTTTMfTJLu9MiS/mP9V64xDEXDkJY7N2+JYOeLE78lY
WvpFKXZ8kYVnC11jaGhBEFdBegfbLxS/Bxg8xJcyGPu21mPGEjaUw8nm3Zb31xBg
bI9FVEG/QyXvaEWURv39rAlAQvJ1ddCsa6EKtsOHiTte4D9H2vewcgT9CecB3GSY
twKPgwgaok6WPVzHLEeIazG7qiXG3Mpu3n4vzLgvJBt8iCqcL58CTpBwAp34z6GW
fbTkj+67z95M8UjAI7DaI2dYcJPXMzomZ8FBdo1RlzIfTFoT5hNllrifD40dF2pJ
ty6ofcgY+uNwUfl6FJPvYTHBO+fEJDVOyJxkg+okS/uCmYP5uSnunuxXpWQOmG3x
+0nvqv8SGfV8RdCH6SVM4ZOvLinPNs1CbImhZmLaBgnAKkMJ69cXzyyF76gds48e
39x3A7+M99r1r/Sz/fmeUqrckGqiXXVaSPeoiMcdc4hE9B/M47UuFbqTYBS1WNL1
yhkIDqiVHHKWuu1zvSGzg/F8YPQ8BzvlQCrlpU5fqOxmpuOM9QhMwZlFAPWZkO5d
j9Mc3M5d9ys9CPRhfrs7ANlR2Xo3jeWKF5GtZGfJusDilYCCQUmBpCsAHaK4XGKq
XQjMATJTCDl2U0J7HXQgXZbHknNHfUA8TWjZ+S1bTCXyxynx0oHIwf+QWSJ1w7fP
RcTLW4lU3jUpwrOACUyb9rqR43fNBacKO4frEGLCG/GX14qvpApun8jsmmcy29qU
suTo4G2C4QlMAy9gMFMBoR6jkVv9PuQboWpmZ5+hRlXwl5+Hh7+3cy+lZYBnMOaN
WKoXxp2LqgkMxtxuBcuo+yyZpTFYqjajFqqTDDSxu4cjAgSFhdi/MLyatZN9hPzs
0cu4cVzLUoenLFk/7Yduab40mEEWzeZmuBiBSnNAOlyKzt+GLTp2YYG7s/IuSUB5
u5LNMEQdZT3jHnlmvUCxK1MFRFb8eZcf7knVwYUZHc8+Xs+DbkV6UndjaFuBbLNB
Jidur6YIGxUpUZ4GArEDMb222gt/c51nG62MrPu3RxOtNRR9byQGtejcohbDScPj
064JJ0BfgLWXAejDEK8DKLZ8qx5RNE7urH2s+EmeUI/sSL/1wEOW5tOxqDR3+pEY
RhwhaFUTP5hufL5yWtOAlxfueO5cLGtd5ePNNjqejUlZmCnyQabfmk/fHth9MArh
HEu5Y//kpWfVAVOkba6X8isMrGQTSKEFrLIzzzwCO0mjkk2ey4xERIY6gzvlNxTx
0TZILB2r71CuPE28zg9R2yvXKmJidnp43AXg+0/bEgTYJUo/GUqsOoK+ngjvbE0B
++GkCKkNX+QoQUqi9ykbQCYW0i7gLR0AIwrkCsZ2BPs3dJxWk2BxcotI0tpJ03E1
IgPVL8ug4xPiX1VKVWoqgTcuH6JwZGODdpNtbg0Pg4nt4GhdHJhTtWvBLU6LjZ/j
LRGhkkL0xgA+1aWJNTqyWEp388vLbi8Y2RK9UsJC0H3zUvCyWrUC8117QNuREWJs
8UgNLMa8BwHIilm3uNfAnmbatjm1WWwGvXYoTV1XNDFZOiODFJz4AFxbx8upGqst
9MBj6I21LLnKk4vVAyQwusXgW/j/QOyC1/FkysoKF/dt2NlONU/Ram7Nb2yIxVdj
URMWoz3xJSwND3SR/+ymcu0tR7Ax9OybzII2C/HJ3LzVj0lIb9XhEmiqLb6Ums5g
m6wV1PGuEvf6Ljq+g07/5TQ5NKX+QeFOwSXVKXAie0ZHXORI59CY+IqGrGSLsat1
JuyJ+3/bNHU/el0ivJ7nvcBXNpx5aZlKf8HJD0zpiHxgg/4ogNxZ97TdcH1eOhWa
2sh2zOthG9Aq6MnOq6PftWqyle6CKcLxY6prZScqF7lbk+/mN/gBjfKKZLTdjEJz
TLlv/qrfZM0vr4uXCakuky6ZMgLaC2sgsnItY/3oT5CNK4ZxdSr9WYnTFcDrNa++
8UjlfGJv1ljmAylWNcPfIlQ1ThluhRNTCu62QkfcEVb2GEBfVo0uuVBt0E3qsIVf
zDJz87Ps7GpjQruGjiQMiBMLfUNH34ELsb9xHiS18729d2U797qxenyoeEGO+wcU
f1c9U6Wn1qxowpmB7R0YKQSP8Ggp8jVQVQDHRUnjNJz4LZtdPg3woqiwwo9BPIWn
tyMbry6++7KeP1g2h9c1wlBXI53NeNiTFbDKmvzRWdCjSCYWUTmK41Zi2cgVzeLB
iOkBjOLjW+Rq/dIdst8gV8EbX1mUyCeMJD63rvmaemKk6kyPUG1HhiwATe1mLgso
Zvl2pDgj0pkZ6Z+OOxVzBzsRoJj1SnGqP80lAXEN2sxYCDMTxj3xhM8RgV3khHAL
4qMBS4cQLp5yduQDVIulRIFJoMGY9ENG6ZYLNdorF0P/JQYAwa5Rb1ifEhO/n9Nd
XqsH32XiPEWoXz+bQ72cC2JQynbQ08teLkSscXRinyIJ2FnsWqF8T07BZt3Uvmbu
XLZimQCp7jbmdiNt+ZCWLrX3TuRUjm7IennAnci8l0/gQMnyOmHR4MGce0qBUpqR
9jv9c37SRjPDNvMyRhO9RRt3sYEXel3cQIKl+eIHWZb/zPyq6mFTQTcTFX2G9RbI
3Qt5uxDNtUAW/8WqhhJQvpuHEvJpJ4EmBWP0xIQ77AiP0Fha1TkrlsK/jpPgYZj5
9/tAprP+O3NHZruoVOBDO6y8BQOWQWuKsVjnktTCpvhefW2jzOGh8hdkSWF94F/U
wljpYNydL84Oeig0NwigUeOzvubcwxiYMXCt9mr27EsS5r4nAkhGDK4Fv8+GHtyg
Ar7KsWukUxrqcSsqv7qal5tD1FbVYvj2GQ+f3FhkhTJCdybYg3loNvh/AP5FggsW
IiEX++F2vqoVePaTFYEECYk9kGB78oqOmZej677FOmLUHQmC7FdI9aDoLjpVv3IK
NBBUIddJcm2qoEs4mGRS1di1xt/ctDuumZXpdGaW2hQCTAAZLFBQXkfGw0GE6m4l
c9grcxnKUObWT71gIXugjMaL7NDR8PrRmualP4vkRJZBS4rPOvuG2oAU0T8gvBXi
7ZnRNuuo9maKPDGinVR/em20r43WKWSxTfWgVxRuAOQRMKmoE5pt54HqhJPLUiph
hPArWGTpx3vrur+9/gZC41PDEs6u/8zy9+qXPjuckkXBu4sNtnaPYd3tBmpbawcQ
Zpwo59RbgYRGQlZYf6ZpunBz5Y0LImzQ6ZQi23EcdNWdgnud1NacG++8DWvC489l
aqLqIq6X03YfOXgmg8qUDNoNmi5xY4zbUKwQLh58PyscefTLdhgSfEBmWMLTAvIC
3aXCxN5JzNpg/8KC9Q7xvA==
`pragma protect end_protected
