// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:59 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Cvuf4KFg9IDJgixEg9O13/C63KAgflDWdSVv+vDEVYyHpyvdZf1WDHfaIxdR695W
aDGxCPR0tr+H1v3EG/ull5gdlAG7PCKIqoPK/BBy9V8y4xy5taGObXi5EZp5CkEM
Q/gWA9ScWOBCi5Vg/SwKf1sO5snoymeBrfTA0Uemgdw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16976)
qd8GxAdbjnYO5CIFoOlVg+ui4bCzAqTw3wT2FeIcpCP23ep926eKxrttpvJKkhAt
NqQgmxmAy+ikt+LLOLWvjx87ifBERLu8RUJ34qw0cS49hIGlEsBUvawNAsHZRQj8
uacYLxl3WPRtVrREB0rh+K5iNd003Cb4e6sGr06O6BvOrZ/BQXJTBjDfLhVJ0jUB
l0DsL7Ywy6RYgIspqiZhtGQmf/Iq4/UY7TGFwPPE2HWTiclFTQLIkOYwkfzqrTBF
QIj1JzKEJcu4je/djKKOTN4chRdeVIE1hk6gHDEZtx3BwXk2hPKrCDYdkR1sTVCG
ZC9flG7xrTYEpMKd6ZikyzGgwoZbI8TemuwXNxMFSkmj7J0A92EZM8jZqyzbCYMT
OpS86tSQ7VpM5Ch8tHGVS6tydME7ERu9F2mghEp58wzBq6CXGc8jxFZnIo05kcWY
KrFHDBIBL+L9rBGZxLogtwPXOX4cKwdwW0ZxvPsPFNikBRBjPFZb7Ht4Gh1z5BWw
IGu+7JTHxZrWzDUnjYjtWmIWY/j+xL7V2kBPXerhvTZf/yiP3oKNmCxuaPrw0Msv
CQ83zP+318l8sQK2xDCo8jIBG2n4hRut1dLvYD3ZFOro7DcGtXktubTK3I/gjQCR
ePDBUmat6TkFcZoqsyREzlv/MvJkfOnEcE4EPsypoyDa6/McCAzc93B0xn5FKv+S
HL3NvRryKpZYF0TnZgdDOOdm4C2KBfxBPKTIRWS5e5iZKNJfEXSCBZ1qNU/hPfQo
8a97e51bF8WjIrmpUfWH0c2t21yEA2bs1ZlSHTjS17V95aPaO1OS2QS3PzpBzELb
cjFxmspSKfm7xVWyHJp312V0utqpAMvtiPR+vWSYHLqqZ+UxrSjHKVagO2hASEQT
R9aB7I075J2px/xb2UFYvcdlQ4CORgRoMuSafww2cJBpxHG2ufs3zchHIT6nK1ll
yEg1uxc4F6DSXq1zMWdb5T4Glbj+8O8yDZukQ6trI5R86ag8HzYBG+mPMMSsvBhu
NSFLx7UcIhlLG5ujLmF7T17x5QSoT2UBhSHRlpDWQCfOMOKiYWZXFrY/d33PrgPs
T/Pe+bo110poXgjxgSzd3OCZU/W0J1e6dxw3kyCcAs9rkRpUcKZgcBGOZ+YUnUBG
gF/h+FanIc0z70onPNp3T614xWJXeOEgJ8ihjsSdN1Gto1gIvfs9SrurYQvmSE9j
o2xuCpJ0J1rkXujtIJNb+A2L5Q5RsfIxDaF4DwubnCpauUU/RhRV0uyXP32Vho7Z
VOOWrGOAy4T+hearHL2/mxiXGLE0kihe/laFULbzEeDkIsSD5mYY6sRFugNuHpOQ
gBn2YB586u7M6L1NvXQlP5/yHwq8vccZVnINQRq4TK1558Wkbta3WVeD7nakG9UP
NJnyRuWJh4QcPAIlTHVPreuXLAMze1VNmY/d1V7DSmdppCHj8S1r7POdvEaCltEy
barAWyhZ4ufcGJOmTorwe/fVJLFY9f93gcJZ2pyYAWo8cnEKW9Qvm0BpFRlQsCAX
s5ShwPqmY6tWcCD60RbnhcnKRQquQVbqGNVNI1VMOX2n4gT9msmfqbVgWhttJT/I
u7p/HWJJOvg5BZG8HeIz3ZmirrvVgMGGjMBwtxfMfnWxjSBr3s/ULC8Bp5n775tJ
0hYy8jPzNoliSr4uxrOeEHIXupcYluA4Ex+DEe3tQjakig9FNpBUZILk763jFxZ0
eXq6hk1sSg6/WDSFZmQactPSfMz903m06kM5bDDDUXZlCG35GBtZZrGn4/YXU7UG
NI1M7D+h5Vbb+OAKaughODj0fCexyGNMcQMIDI/DdWfZjtRm/d8RsdDuBxdKZ1fl
J22i9hW0VK+diH3pPErvPJM+O7j/GW9yynAJetlbi4fR3e2M+7OxxX8b201MNLr6
cx4DxVZFna7bgcRsCwEiCtDd32KZDBxrbKfPm2TRXFQcIXgsBuegmvmuaJXuaPVm
8f7f4+BHYTUZvFcyRRxba/Ek0BX807QCcEGXNHgX5yn6vNlcS4r6dN9MYg4BfmaA
DwD3oBdJi0QF7YMY4zssZTyZkWodquVYmccsWgI0O87TRMY1DOjoAujjEtcTE6Nh
hrkvOFjODSG/b7hCUWbYHnRB4++XU4EPbzQtpN2IU1p69FeQdMwxHmpdIxMW9Rek
AmoI23vfBpYYSdRPaMLcWa1H77Qt0ldDCx3YzyeFX6wAKmDXFXzJyq5XGFyJmrtN
OIlxgsozUDcPEDfR6Ydw3entmtzC2PMJgMp3+Je0MTgD3/p/daapDnusECuaJnix
D3XB3aArCFAU+4rPS++9sAf9IP773XmYyGu/t4FmI8VmbB7ER5YoAHFhffxqifed
xbAKLSxV2dlLySr2SUbPR3IuaAidIAQMRRehXQ4WKXZZxObkQMEEukFa/ALh/eQ0
wjq90x7GLc//ZkA9rV4aIRhtVY51QALn9DZc383pLGGvOxVX2041SwFYI8Eahrsb
NHm0NiaWS7M6uYSirECaAJFnf19pWLGM++wZVnXOIdvkJ1uAgEGo+aA/ZyAWg3MY
mIDNx//IjhLjSNWcLUllgV6gp86l3if81VZGPpFGW3BnFKZZvcRqsC2U1oehyz/T
GtpxYhG9s8I3P9gRAhIQJUgzxHIpPMN9N3dusx3XmCwvKvoEiknn8AXQ8PfXi1oA
UcJemMVPixtX8lPQTFiuLqqByo91xEX74f9u51aidCCqRnow1Szae39OSKjxMcVS
7NffeyJUq5vcnLebYg0l6c3rZZloVy4ypfvIdzTHZtYwZJlLw28nmcrXxG00JTWc
enx/VVyXNNfX2CZUtXmDYTZ7AsADPEkyU2o+Jm6scgwIuHIHA4siYn1DxFQwzo91
KxMt09ZH+vYKr11AFMuQaWMmxuY1GcbI9WfFngcAYUdmm7Khk5LQO+WBbRO/ZtLj
0QhTZLJ+G5/8PxMa6nMcznj/rPDJ1jsM0S+J7p4VPkuxTrSMrNJn5gBGpFT+g3eU
Qr7dLyl1adM2C7AzZthhCybQRVD4KvY6L4VYtRKkgV0J/NPTZvH996XXpbWeDsR8
nYL7Q5VaglatqVVeX5KYiYL9OYuUMKl3cKNIGpe5Qacsdgr9sEK48KecxaIhcI+9
/VmNlYwbIyRQ36QRaE0Xb18qqWFBBnSPgjeabF7b86Wr9z21hxLCBzuRUwYovF76
ITC0ZTLHM1I+RW9npnWaudhdsHVScsp9BHq4L5YVUwhu14VhMyDDbZY2fYCYEyk6
YlpBFHn1gL4yHgmCHzmh4jUMP1DhHH38pAd44RJH3hwQl19kNo0P8ilccn1J7dos
Qpx2MnLXaknO4FOlgivVUeXjKivw2uYCYU3O2V1tneg3UjvtyZPdBqFCl1KKEW3Z
bD/JhLBsYDC7jFfdekvJK6aStlsGg+YPrjAe/H7BGARKfOIl/drlfv9Vh1+0Y+D3
kuuzMmAXDcEaVGt3UBiTTVXgqKLJJbJnKJbh9c2MFhQA+gpvW/GizjAPPpUkkRdE
Up4/5YQuA1kqGAz87LIcmvH9SK8dC6050gbgFtccD93HaCd28vccuIcfwvJVUvfC
QFVTqghzNRF38ZTuuGEDPMovRDpjY9iP1uFltSDzLk6tMqXwapg/lYXGxeAGPKUi
8eyL6B/nwBaciE3gFuF+7UHKHqUP6H8mDMwTzseyM3uxXeaQUcuRSSJ5Dh7OwPTU
eVpNJ5Tolw4vWX1d8awzu7Ls5ntb3o2vsbXfj9Q/F7GLnKLvpIQDQVpeDnuuoeua
Lxk4xEfOsCrN1uxY/FAlwBHGu6GtdSzNjFh9MddUF02qcHl5ljzecbWO0zXnlnFc
NcVHUBEWKaaW200qRY8mrVlj1lxXMwXVNGl0cKk4VpYql+oId7TuvK+KHyOP5r2/
nmMVCpTPe8l602YMBmxUM6C1DrO2C5ksKoRNlX12DQWS7s5jUycxzPfY8/R8ADYV
uJRCf3BFT1nSCdRuWh81Y2tvWjMmmz2IZPoATfaJqiZzw5uGupkb9dJMkEq36Nub
HR9v0geYdgABPLAoMP4WjXf2jbT8hvTXFR9AIs/Qkoq6BtBSCVRq4zDdkJraG+wG
35GW2LwZCyRz5FO7LNeTANPb1kYFahxwNUA8GfUMyv5+ZJoMkU1dLCRf4LtBB3QE
nbGtC6s8NbHnY2SD+yNb/HAu35NJCy/edo8CN7i7p4Ep4aiTTXsPInNXzV0U07SR
yBzB/PHRJVUkZzLIGErYSkSMlfS98mIKEJv5YF2f1db/MnbB3uBWCvSIb3ayU5fN
JF6kbM3AMEHM8jLgtXkkW7bhxgCuEDpfb1DIvMBJjJbejJ7Ph5pU4MlnI1lDA7OD
sN+TMbVs2Z4iuxL8dgzm8Qm45w9cgkHmB1iGicbUs/Tq/SyC1E5lIt+HogKfUMCP
Ni4EqJzl4TmqpbV6XmZUWjr6WncvsPPZKHFwVt1CXfFdIZiHzum5ynPX5Dh7zR0z
2/TRT0I9LJhqRgUoHmQ1/B8sury0gbKG8HPTdZ6tXTek9/nWxIVkfliwWH7m3CPc
vnp0txpOPeFrzO4+Cy6o+0YJM89aT0liZ+ihCBedjD5FUrCx2StQm7nO+5GLSVAg
QXk6X4TuEHfhawj7DR4qwv3Ty4VPpCZ8nu1NRc49ImZATwxS7j+dQuwj1cF2GYGM
I8MDE32uEOc/lzvz+Lk5Mhodirn2UgNOLSteppLxOvpEG67lezzMkOqf/9LjTocp
GidfohMQ+fXsNG1dJoExOpI7/Gq/XYF48uVOB2y21dTK+qy1mbAB6J1wQsq5Bpp0
mrXnlMrBt+T8niIjIn9xta3ToFftuk0qayF8eC8DXxWXeuSbnIa0GF7t4iQtqBLN
cC6AaqQRTOfaTEK6avboAo5ezkfj+nfCfSACHlwVpeNJZWxmAMmukGBCpKMtP1XL
G5UAk0Aziy/zqQpGutR0q8ZY+qdBPHsBmau9pYnBwqJHAAN7Gu4yzefObl7+QsuC
Vx7UPs4WfNEFr4/fvTdiflsG2UlAwhhKwwPHYa7Zny6Ojg+1wyqXL0G5k1JAp4bs
enuGASJNcqlp2y6ujA/kVTUNgHrtKpCZM5MHAsqUQPRLBcaBh3JbRX9vGXqO/U4k
OgParBosuNB2hGu9+/3HGpg5TtGoLw5UbrDe7Ateub5u8H8PhfTPVsziOwUnHwMF
elbw5XppKZXaWl+N5DbwchklkM0SownAE/1FGlSUkx5/8g5HXdTbnJvE3T4GvMuf
xdgS40gKU+VCCdkO7XKqf8owEKgSrAYiNhVI3aGtWVIh5TGKjxEHdCnPfNFyt/Wc
sgb0eER+u+GkI2GEY9u6EqgViT1GKes0GeNMvxIn7GSgaerCIpQn3tXFnvvhVUsl
Vs3k5/JzQ+vpcadH/YLqnee1nf7PhXdlyFD1QSmzlpqNuF50YBAQ+EoxpjaG+63u
q2ZihUK3GmH2+vefMgy78OAf4I/EzmqaEv2ATYAZAl4VL1NKG5X2S001c6CbW9L9
bxmmOVYWBs/Thtk6B3yvY3NU2fQD5iJQQBCZ6vK6/FqkxE/ZFfDbrDl64VE2tWs0
vKbm3GaeJZ0FGdGYt3VuDVshMi4o4w8bQWQtbba0iv3iCs9OVou0VcJU39Uf6z6C
lDc54Stva8j9zj5PzgUu/XUkOQ1X+cAfqgyjvvI93C4NPYylQ+nxaPglaGlMqHVX
XdtqvEJ9hcbBTLhbe/oq3tw4GDwmJwrTwPdZF4DJU7W45USfEjURK2EUA93cuYq+
YvGj9KBe8UkNkZp+ScmJ5JNTQp3ncelR+daHzusd+kmp7mPoaPlCx+HFmI+owkmm
nLT5iJOzxi6hJZRmtLyuJtsLstXnpfHeChrud83vmAnI8Wt6Ejimlnl1n0NixGM8
fkNC2cNXwwc+xS5xhtnUzc9GmwbuzPme08gFcchInLP3URyIKpP6n2aojLv/vBsO
JyghBofzFLYKlKYxjFPfKtIDTEqpCqbS0WSKxXMXXzqB5XVL0GH2AQzqC3+m7YzM
2v7W7TYofqtkhYlvuqbVI0vhEzqDwmDed9OxXrsJ0n0kgzkHa4kQ8iq+2HESenAY
bDVniliH7Sw/Z2LoGM6LDJgO9PXUAFLw6X1W2php+UxqVSi9icy63B6zGbhOhoHJ
ztRNN3i1reamXnuCqI+b75mhKvfogHOyyprG9tZbxX2KbXVzah08hJJCpW95HxgY
BWFzikYQmHYJ2NHckTiFrE2EQ773w4B7aPE0C6yQ5O3n8QtTsaqLEQntunZXAIcp
IVF49vrvXCVsrbLMDTLRZT7G6agEBqddle/15Qc1Dd34tU4PDcb8tb2KfvOD3n1y
r8m6o5cH1SGTk9WVCzajYIEgHv2ynIoiCKpv0AQ7/7J8sWPH4Sm4Rv89ild3fGgU
Sy9WuG+t3XUF/2xIVeXBnct+2+O8iMkw5bdyzg9tGNdXZcZ4ibul1KPs40sqeEaF
hKxqUx7DydHV9JeVzvToKhxOzz8/6xwACX+ftxmJ73Kdu4f0boAbXqx+23r6qou7
83eNDrCn9hjUN3cx9JPSrTCAqX5n3JbFOVKo+kdWoPsQFwc8ov5P71nL2faNLoqd
tKSrPR4LU+T1Njw+Qs5ZGYUWXl4jEWKhYmVrNOsv4A9/PFn/ZEgLyxXhlFFNUHYY
eVtpfW5BbLvO5uKe4b+ky/708OFx+zZB55/yyf4B5rClv98jPS2sMqsObGHKi+BH
2O46nKOW+RU73UNwrsVzGR6UUPsMatdcMpIK9WsP7i26Vtqi4hp7ZFmjBCMX0SSC
nGCo/UHJGN7Z3PUEta/974ggtn+hvHEfNHrAA2aGwtJLUd64F7ZVXhG4y2St+mDs
QOHngOe4kI7y+h6qg8P+06ZpEsLnCzykHz35lO6Wln+GSHyuNkLqiNJ2Nq0xHIa6
LvryqEXcdq5QPrFsDhpfAbz+wJEt2BIFXcuYLIHVzYaerVIPbFB7UJLHoJ/qqCsS
ih7oVXA2hw6xwHqTruMJ/NDgXlI03MTvRCRmoRYPlQ39x5rT5PJnDIF17oTIHlNY
B3et2S3FUV8BLXFipzFlQObWKv/sMjkuvF1y5P1CpCVfCULEfUa98BkiErTamaAV
MlcA8HofFBsu3t+ctquE/oACn+uyyX401laI3KvZ77CAYRs+2qdJj2mefQ8p8fo8
xrdXrzisU0oVBTRqfW4Ya8p7SUx3julUpGVCexRzQqIqSQn5mWbYSWpCNosDoucI
O8XSFbCa1PCmThUiLS/pB6TRq2uuPWKeaUqCuyttNuYm9TinxI3lm8DfXV0Z4bh1
1N79v0XksX2wt75dNha1vwqRe5P7TtnfuMVFZZoyVf5YJuEwyLrymvs59Zae5+0h
5AL1OlbkK+SSB5/vrVpFpbece13KVCssyGoEa0I6zW0osYgqiFQUtJZgsJgPVOXj
STJIy9edzkscYBrhPJt56eabh3PVOBMEs4TUIwyy6xD40tndlxF9RokMH09T0TR1
vOS94AIDWDUqR+tK4bgKZ8Kk+kbMyTKVyZ/jjk5Onu7050FuMT3ID7pVtP0A92tx
YnS2LQ9Y/YggHN1GlFZxtRxeojDix9NQR9cQMB4a04Zn0P4GbPkm619xK4kYrw8i
LF8lsItWt4MvHl51smBdVwJnhq9G3ZBhWwWHWFFQ9YHC3wsOQBYtMXvRlQDcB2nT
J9fpHww/rM/7omJVfsQwwXa1AGVNlqTQTvjso+VE6y4/yzi+1CQmlauYQUsXJl2A
Krh0SFU36f+HsuglyQcgQ+rxocY6cxSix0MW8J7ujR00ijjshK8fSJ5xm2xLEAUh
rxw4/o0NkW9pMKnUvDy/CgJwiQd4HDjF8bC5I2pj9OeiNjJ7RaxQT/xwQZP4zDVM
MLfpRX8HatGoDRz6Q9dW6PllJFfmAkPG+Ryrkb7FM1+4ceOUZyuJGNGCAtuWP4m/
qTk6u/bw/EV/xxLvhjvKQ+ylVVVDVyRwZcMJ8fnTHlTi0rhU0bzrtu1DJUyu4yoA
mf/CblB3uBa/VUg1J7+cBinsgk+cWoBBZiroywKOXlfzK8TYcN+jJ3FcpSNa9ml6
x9SOXW4VhquSzVXMRDlz4j1/BpK/tZVaAwyIqOUODKgVzecj/O1oHHh8U8s9+xyF
eEQVbbA280oU1WgaZn0Z7vfO7BqELpIMqL3LHxemoYLzcYUDhJsu7a9PUhu9mIYk
owaCol5HnqM00P1aY7Ndqcj3NEz3gp70cNyV+VozTAzjMkmV8nr8LBDRsPDd65Ta
D2aou+1ibiolKwO593tVHqG45Sg5iHe/OmQQOrD0al9QTNEnGk91x9UT1yTEWEn+
/Sjfomhq2yzfcUTgE1kv4Hgo4+f4XYH1aVHVzN81yK9LqnqDHxjiMEfQR6UHw8sU
mUNjs50sUznKAucCVw3WIcZZfGlMQufgfwgVkRZ2mWF9EnPzo272cHSmC1Q0ZIGa
Jdg6MaU6SYeVv7IycZsnWYpCrmgKx7cfKdUGqtv/oNnerBICRwXHUkgCPl/noYfv
MGqWsLC5AT+WgzxW0j19Do2Fx7OVd4mU9yOXsGruwzREUZo8TG6w8mSEOtPfU+TD
DjR8m4+BaYNjnA1q/aRh4GVZ5jKvt/XZ1FoaQYkg7OvxKQDByoTeYuoY7fVQZ0Ll
zljvFSjUc7/vGwhK1AumyQgiBU8SiBr6MUhG+FIG+IguJ6oQBxJvQcA5bfSQfptp
f4e9eLYpRTeSuWt8r/k3/iXJ0F4cWTFPoFgiuVxaq7F8s4uXzEaWYezHWQgjjHxu
isWL+BO4VuYFAC5QINY1sSkbgtDq6IjDuhi/nT1qH27ivwFOKkxEI9HP616Goj8S
+o4iwLS7SWTtiqxjxgJM3qMkRj6N4skyhGHNrOL04EazR14nY10STUp1dU1mpvxP
jrzHJCzJN1KJ1iAgk/DegBq3bo0STJ3nTam6mLpwcQfm6lDw+bSc/unQjvr5CksF
SYNgWIKUgYx/jQVkazFkROOViw87+SeEI9FOP1eymngY6B3i5RnR0mSCagTtVmAD
dAJwEWEQ/mJhKa5CgGmJhAqObGGkZ7q33XTn5DTtWexMVsRhU9iKdiLDYtG/iy25
Bw01seY9pAjM16yGZ9tCbFINgRa1gsYaPzr47AZukSmNBAo10I0OT+6bqVWmEx9f
/Zb8T5W9fP7dP+XhHYd3chu+wIL0NBV1qOacJz1h55BpVbqdFGh77/s4Tm/D+Dtk
jvU4OpQKljOjIc/yyf7aVkokf8jh3+BvKpAzAt8xj3wfuSefsUn+DYJBf6rgZCjz
FXLsrZzK9gfnwP0kB9zhk5gMxphHCB7MNpBgmMVNtHIK/2q2W+Wtgnqg/RvN/fVm
d45j5WlYor1bs3arplminzK841cXPxn7iR089SEdW89qPXlGjpNokJ1yVy9Ew4oz
aAJHx4AfVicVWaIUCwLqkZ5ptYb8/oeE06KP7NyIMpjh7z5n1JOa/GZ/d5L5DUcs
C0qxcagP+tQUoLMgzBSXYeVoLZv4QshlQV+hhlYZwMH7WaPgsyiRRK9yA/wp8Wxd
1KWnMur1HvcmnEwYbxlvMMiEVHCzTOPr5DiwCbYkzPS+FeLbf6MR6QV64ARqTcnj
FLPxG9vA+NMWAeLDwd92yk0EiiNdVqHLv8RFCSjpwDGqjz4lzevJdHknhss8Dpah
8y9Wjd+uY3DgA1dKjhju/7xKRnSgt+BjD91D5RctWXwWgExFNUPtZm0Z2xcY+rs9
9taQN6VAEmX/q/eb+DHFg8W3wziKTCm56P3ZQsgllf44uIAWuRnwRjntua+/aRW+
slUOsW6Mtk9ZiOTJCNJpAOcQsTDYvemNKdAZP9BZ9VP2/GSVMT2HMPFi+gKBvtLp
Gp9nGe/3FzNz7X8+EP1IW/ViV6Rx708tK93oKJ4kFILVHVk9Cp+3a0KkPg6wOH5G
gSV6VkBEvei8l2Z6acPK4ZMY4d/k9czsa0psnIJObj+eEE6SUut8VXXaRMxP4bh+
BmrUQmMQ0dJY3r5rAihFrp/YEKgBLfHDVk+qwkIFKlx0nL5/Tv2B/jrWDrlSA8Dl
M7UTwo04LZ/BmY0ghkcmVGMkhNAVtsY1e8fzF8roSX410iEBvkjArm+bAiBD+O+K
EiBww7q17Ze09ZvI3xbRAxURYh7xhfd9mOxpD89NWLxYL5sQWJhjOZdt5fNqFe58
GWQvZs+1XLoIYPw1YodkHoQrYN5BbF+SKWm9Us1pBKJRw1MCNaDN0yJvVotTPmhb
mp7FC/45phOHtcsnXqHmqpKLLzEnd5JTawER1ZgMiOSkzwbJeOujV5qzBxLvCDxs
wSjjBE8g0hJFYmKgcQi3koE6NVfz+UohmQBwbhGFkwHtjMolsh0b5lsK1queg6Pr
1S632aKBIEkW949F80Bz1k8GNS7kzvLRw4SRuN/RUcWKl0zf6tOQ2DRYYxpyhBBb
Oad8F2X1GJHgO0/6dPp6Z9p2Xg4W5497fctzVUBSsZtGokjqP15Q8CeICEE89bvm
7Browlk1++rn2ZFWMJ32G/ZWoR6aqeYSbY2KiUdPviKz5lF9Q39k0q3L0/8wFiFV
15k7ABqCC8hdaHcX2CqHr7c+WHbeM0NdNZOvbO7AnThgQ38+2xX/hI0H5BGhjssn
vNlHgVgbM6RthvnLWN9wdiORVD0ENaqHmbhZx0ApMKO4XueGJP6cs5a2LQDBpquB
R5yNvzQwSkte1yRxMZXOItG417kAIxY267SOSW8/TZaOrlbWX5/RV1Hh+UC4nzyt
I91MuuptNM0U1dJTcFoMur2tQRFfd1fDKWso1pgmbwsv/QZwv5L2aK0WhkHhgpbi
qymCWdCfX0f002RWwtk02+ESASxBQIBWkYIB8qGtkeTA7Rwo13k/BBBU3EysiH7b
oDqHHDEBtQ3sAjDc4V3RdtuF629Up7olziYIMEBs/24BzP6/y225LM2i71Lg5Xvi
8ae+JG3ik3WgqMMPEmwAvi73K6Wu20+7RNOryVRu6Fu39vQfFRzamwY6EnuSwR7X
WedxTRc64TAwUOczziKkjdPcuqREK5koVpy4uPb7D3xcDe+dcv9H97B0T6Ab8dQK
nhoIlLODczond+E5xklSv7XkTIuyYdACJSsQLGaWggK2SY4c4xlXHhvbTEEFKPfq
oCSdeh7jGKrPP6tLmLIVreYSsqUTuN7m82XPPIWb2LQhsZ8RCygGfInfeQ0mRY2w
uHBQb9OC/N6tYHDfXJUdWLV3KDCSSGgX5w0iELEJTlpoRxe3qJQ0GKbdzwLrxLLx
cFK0txoRG+vrJ3jQ5eTtFIrVgSCdB9ISs2Hx9yFpQN8nq73yPh4xSbE91D1F7ZLu
7GkoWNs8STJz6K+a9hATzZIM9fuRyTeCN/6HQYbIT68DMY6/CO6YqfZX4FxQjgUc
vlgn9KFxHYKfDD0m42ZI4OT+oxQmFbQtoXJ6L/sqzRkyYaAFUJDVnXpY9YElt4aH
5wHLULTvbApHZikP3yEMGVH7mJ7Th5D13X7XuJL7spSy2r+QPrpnIVF4xxgW9XkW
zX7gehfUlcf1wUGL/4HwtHqGfQw399QkKmNW74ivLu9dJkG4CFDCIdV6WK6u6CcB
5k4xaYeRilS1WOC9Ku78Ub/GEf7HwxLicRB2LnwKBZdEjTuw9NcWB9Aft7OBWAbX
L96/KZvAIK4O7H3nEvRktr6jcW6VOq3PuuifjLn0L3p13hqU/s+WVkc6RIR/ZDAG
o/gt/pVynPGpqTFJ0NYOZ9FErUzIHRcg0NLHtJ9ehd4CNsKYTHGOh1sQiGP/xg6q
3rWBEMX6B8glisK0qCRozfxIdoTUNNM6awHvwAoRg3/2x1GCZ4zUKCztfihATfO1
KJKFxfZ/rtvFnnmFpY0/pGi0XPfDqbEa/85ZS1bd6gXlEJiulHGknvUJzm5m0Jss
aitxxof+Qt1+K3OkWuZDJ+6B5y/QRjKqC4SzzgsCCuaua9WlHSMk3edLnU94YJwg
xXzYFl8FrWZTHqpjpO1HB5yR72PNucwetadVcD3JRYFaJYoPT3HsEGeH3tFv8oV2
nZkZmlwHsiBw7kqbOJSHrJC9WPSgiz5zmjaAzWr58n1+YHxuzPcKRDAnQ5wS35xI
3Lk93j/Aqz4muYzhIspPJK6HRY8wrL/D0XR6/I6S4YZeM0snxJfY2vP3ojUQkuVk
P2nhBxHmljEwAEPR0OJ/xkS77nP7AM1xLfe4dVXsTNJLkOun0m9APBNse9ZQ99hP
Obv1CzzwOJQNJKBZ8YYAOlIbFk7i2lGGs9qmdYRM9/BDsKSe10pQ5bzFLb4PKXXO
2L7XYCcKmqxTh//op1o4e/C6InG5mVZozuv3LhNF/+OBBoFeGLtQDK6fwikpCAmN
hnVggk7qQsZHeoh46v/HlVsM6rumPEFfKvi2d9rpOFkmVPrie8xTg92rWqj0EED4
LATHFoIeq2YmlRf7HpAdDtyOjdpf8lqdd1AaoteDvrs11bZuqGPIBY9ORPV4QF2b
iZ28Vqc5Vrkc5ie77GfPnnrjxoQgsvmAI+6stoCKUNWW36P2r1gX/NXGiPlUyXlH
Ph7HM7uprkZGN4pYzfoaFFeg+K9IdXTppTn2/QHCmEYPfkvh/8pqcD/M93Wr18BE
w89SNkqZZOAYuF866EAcUresHZI7nKM+AHkcYJV94+dM/YU55iKjZC31opKulmAR
bCOpVCLPBY1gj8iwOkhAiEhG0Vt1lc5ItBo86u2CZN7ARWx/x4Cmrt0l3NzcHSAN
zMiVWg0kPE9MeFCrWxn0UZX8jYE4OyclA0ui9Kcp4bnDjV/OTDbtg3sPrS4rrNYy
Fqs18zvvjBn1kHT6N39e2K1rTWo53cu4hUIQXeYCqcaIz2kA00GapNpyETT63tjr
TaHEoa4Qa/glBrujIfCf4OJixhovysfZQUG9oe5Sgtq2LK6OD2TL826AtV6dUAUS
kXi71E1yg2FOKU7Vkvin2uj4fELypIuYBkCGD43FcH+qDJv4uumkDTj38LgW1Q7n
IPfKdJID7A+XCDUpgzi1QXO06Dwui/Ur7H3qElDxHCQA4nu0FbDfeyCqFivYcUYQ
ISgln+ozvtnDVGYsopXTPzXN/Qj3menoViytzmor6ZSFd+WTy4JI8+Ul2jBodnD2
XJMcURzQO4HhZQcsN96RTEJRxN6OFF4H1wIh12N9i2+aNusTM3pZg8/YzzTrslXi
/3vCSAkgnoeNuAWebEfJi+FRbohDUp27r/bKBviVmAH4brNVQRCFEqeJJ+z1EjeQ
KVIbVu5vMDpz2mRqJenr09GIgd1J5s7g+fwXVWxRW7S54pLBxulzU8nme04DXWqU
7FuZFbwHVcgLHNAkYWie/HFpBHqxo0+D4ChVjuLZ5k0lGMrxvMG2w28ApAnCsgHB
BDQNEah+0KwDXEkh6fG3ZBSCWFAzkS8xH4OCj6LJ8hwcz27EfI5wzCTSWppDo75N
+nck8y6OlWGy5rCq941vwjFbAqcy5KlcCrD52Go+J77pdPvgqvdn1uH9r5tA6yqD
SPeWGAmHCY+ZqF940a+lKsTZMdFGEHDsqPYKspnbFIBGRzNXWnpn1VZO0dxrya+C
m0hlGyq8HLJKk4Pb6lAayn9BekrjZZJz9+S9mqjlIVDZI80sGtSZ8bqCUiytGmfN
ffX/+ciVADFmqT2Ck0nJ/RaNJ4YSM0G9Su0Dpt1wkh9XKxLkevPRA67xI5+Iv/Vk
iHmtTalvbENbEf66MepBcl0oA4ez/6ON9xjK83Z8BOcUU9KMvSlDy6PlXoxiE5FZ
C1qK+1lfBYH4IhjwJhxY/lhxSwPi8AA0xQlyZnZuPnXiTlOdLYDOU9UBzbFbt8aR
kVCvI0RKFh13XDxESZkAaWM4dyyRLKw6Y5NlqGdhTLkP+wHfBRlwH7CmsSBEtRcI
/zBGGgPGLgTMfFZHaQiUsoaApbtabw77bxGOulXRg+d1hMdE0723KNyf52xJ7KTq
20Zubu/HfLMtYc7mu6GZxbHKgS7fIT4lvjoO7wyU8TRWrfulcK+s+3dcCAz6gusX
sgTQ4hpn0gcM4jMUF4puCOJoC8dHcDpximrLgalVQNa9GjiA05ueUnrGv5IG8XvM
dvZaGIvSol1A9Z/wszgYlt0+S/0aKk0urCvw2QpyHvDpkkHrE1yd2vn7HZgGsBul
dorKCmG5n8OPakAbWL/ImMlV/1T3wRkN72z0iogCMc07kVZrIssPINyXXQfkhxGv
vhzOHTHQkSIMtry4+7EtKKe0icm0tIZLwisuxfYwOSDbJIrnhX/kvnn4FOFx6Uf2
f44fnkbSrxL/OIz7BLFdOapOSh1xU/J7bnszSDGPS2MouKTYPRyDcCZqsZNE4Izs
cpMvo4TTLGJ0TEcLHiisHHEyW78lXG/1JdxDoQ5eEfuERpBUJLdRf977IjjqTWKF
eb79arO7lMhuwgzqZ0wh7f2e4kuDenSh6pN5Z9+p2D4lJwxxeiowylNBFVi8YL4P
KNl7WQ8blSUGH/p3j0Meh7dA09NaYkJCa5H/eL3Rw3DV/MRIc3jZ5EISPLiG2toJ
UtRdhUvueKvX5bE2J5UpN/LYp/X5VNJk7NIt+GT7A7L2n7iIoXQxBiwm3XTKdybv
zex53LE8Ng9iLj8SFRrfNAHH1YF2BGxawU9zTKH9crdMM4wRdQuPhCY0gboiNgJz
k1W8gVSH4iMtoEVVgNyieQHc9XOdMpHh80F/DpGqnkCTARB8tn0nlYk6CD1Da3QD
ZbF0W3MdKT/IWIxRA/eIOJtXX95LMrVdQ/Bzi7Kiy/3S7BnjCHhseEDFQwGph3B9
+PtGwk2TdEvCKtZlm7LZQQy4Se73AtwtS3HMABDSaRZ8geDzJtHyG+WsgXFj5++z
qYT/DMQT/y7kFDtr5xGfla5Vu3CWVK8E4UNEfBUNxGU775bcBZ0nBSqVygp41wWY
615XZs77VVB1pfVSJP/8DDqzt0S4ZOnuspA9zljkpLOue8zrVJWJANhyQIl42ppR
Zbr96zXT+dHCFCfCX459cD8iHf/URO+/Akh+IU+sVKVsUZslMYXnQxefJdrdXEE9
v++j4ydp+8oJ9g03tKw7xfeXoNGmxYcAHClTQqZkJI1mweJ3ahnwxgSibAjtLqqw
sV3SzcnhROS5USxyQUkyNxi+gLsxrLnSE2EGv3e85bbszQ7cbTj2vi7w7+mjSUR4
7fDF+hPbvf5lhNAiK8tk2I7lHK52lHWhETQXt7xEEw23PUnECPz2EwzYhwA/s0il
Y7aT45sItRRDup50B/ru4j/rBBSRVh3gYCnQYgKqq3TrRR0HFZD4HNWhn9Ux9GQu
Icd7pcNhM2w9Lc6mxjylLitt+j8smiKnwSo4X4Js479TAe4KCGdJ3svPLOTEZceZ
ohc9FxMdxQ+qh4BTk/dpoy77JsvSdw9ZR2d4aPY4d8nmYlN8lJ8rJMnjBTqbkcXg
5Nblk/BLgKsUYVQ2JIqWfQQkpJtmvIDCplJZKOjXAO4MT426+9O1UV1cF135owaN
rg+xCUELrkrMYjPCiHgAyU+iEVDjsg5sS/eJWL3VkkAoyK/9OEml2TUQD9tlErsR
e79yR4UbLb+jH2ZOlhsLw612mQQHgv1ZE3aRTM/PEDO9mlEDb3q9iHFWJRhI8rHU
fkLOfoJbJAQySsz/rGYx5wsraV6+rpeGxv1ejkvY1qGqub3YHXqKtsZp31sOMZO7
M3OmJromwVdhARkYH5Mu/sszii09J6XB8Ln4jxXeJYFhAgiNbgXpgbLKta3jHR1P
X+EIld+2KEQssP8PG1dZUE2k2lTlqSqdDArH1SjKu1i21MrL/dwjx3U//WraT5Ra
a6I31n0XOdo2Fx//KWeq5m2e3Y4xJrA6iCoNEKpqiXw7RCry2zyrYBSWt5tOyrX7
a7/CRuyu2teWcoZhYCXfOUp4kSXPbBc+Hu98X8Gcp/irkPLTWCsCI4Z5fjeavUNb
gJKHvOCFvOP90p1msLsEZ6TlCtO/LT2HxajWJg/7W4ef0WJfXEG+2f6vtSRJwyk2
NZuL/ErkeN/GCs3eUWV4yYkVwGPUeEt0Tzo33igg/qOqiFqKjxsyD6T15xdMO3Mr
NVGVpknvfELNwqcyJaCMTO/8ysC6DmS+ueFHAdrHdjFctqvgXIWopd7No3tZ12Pk
2Lks6haffZxEguHYwFAsO/HGydfzGsxBRQAww85636NEpHHxMt4g37MOI5anu0ET
X2acu3OTNL/I8GaWXSUjAKFd5TiRcEmG4IsKCNoGqUT/Y/DPNpaRunyg/GDb0Znv
9/FmBYENa1CoM+csG857SxBzmMxoHUfBpN/Ax3drYPLmdHbz1Rs8+5gqs9CnrJ7y
ONZtnl3g8I60rWbHf4+PClOBURu9Il3zJgxpJffetLKifIREE/wYzvCVBUUXZtsG
z8gzMQN1WNu3LFeuzaA58HDx6bB+1E63GR1b01sWuoq2AZZmNnGrM0nPTQXs1yRK
lOpqFqCy/gjyqunEZoPz1+aVZDpD/NUFaZJT0cZOFajCVw62p80zYR/1D1cuv+rA
limOrk5jHomKZWe2DfFvW7o3ruCwL/W+ne91p41eUKKN6qV9E725tIq7KTixXllK
ncfUpOpCrFpAwZqdN4m+TqnJ++/UKD9zIlUvitTTVOl4DkMbpZHvuDrSFGrKWAZ2
fM5NKhDRiT2psru3XudbXKXf/km0AJD/93yjwSa7aAYPLVk47p3IF1mkXmMKrO/K
I9vW04wcOhF4RzMBc33ngiQiP7D8Lrg1chNTzhzaA8JLchwIyeOk/EtrxlV8kOsx
i3Bk2GDN4Ul82JY+9jawsWZRKn1Tdl/CqPIqc/qQKoFGtMZOBL/iDFC3vPftMJAe
oxDi8kz9kkbpvL52PXUUdztIwNcaX9zxzsa7X4aGICZVkhqAw/jMviBoVGaV55OW
AMrtG6fKfar4a5hSjXfGTuSJdhOeaFEa6S1N25FbD3kDQnZnwfE4chP0aTgK7Gap
t8F7AQQvCj06+DbcuItfiBZVVtUE+RjquzO0usHN+Spe5Tuf/WniBfRxkUF8m2lU
Q4+8MRwUCWBCxTTgquAj2Mi++nvmf+BMxBjHrPgrv3hlZ5XDb4UCICs7DZ2BY+N7
FWkfUcMKGsclWhr1KWy0EGpy87yRSXfC0e6BnFdGVp2xSATi6Caw8OCNMnLvLMJz
aNGAugpy6QyMsZPJ6b2TlhCQ4+UqAwQbTgLfHixcj0emKKdvNsnaO86rijQ7QFFl
mHJ3z7UoP0QWYSkD0Nsq4HbHHX4awLSbZc9f4C63+d5gdOC5k3PLUYL82Z58qO5E
5vA52CVxTgV6QUJBRyhTlnSaakSvj2bR70psLY3LEYgkHxbviY2a11izxEgTGZYt
BblxEP2Q9liOfgju72EKf8O5jRAsCPFAQELDWAJPLjA7D5O1JnSnTXbfjftFJjpX
sdZI+H5DizDExzIQ5K61xb03BgGZDDTbhIn/wzNyTnv6mwrE4OtLygwN2yuCfj6f
Exz536JscsUS4LAVMKuY8HF8kyMFpS5rUaOsVp8iZFIof7OvjX37gNtA4p5s/Wg5
sOroAdbNkWYQzHT8s6cL7zSQLzo6EueSO1UGpwDiQC/lVC5wUcit3eQ1am5QDsXi
+p6V5PIsJX27CzsKevua1MG8gU6Rc1iUeJpIsWs59gVjJt6d0GZbdo+e4TQDmHCJ
/zqLH/0/u2YaI3f3BX23cH2ze4qwPkmb5qXSw/LcS1PpUmSmGxnzbJPGfCeodqiC
/Ms6V6GE7nLTKJRJurvQ6+ptkXalYDTkJia+vbhiuh+FVCnz7NZL/d8bcbp4697X
76dl6OqFY0agAr1eS4cXhv0MKvzrasnG3uQeWbx4d+ES02D2YlyB3isycCG1mid0
a5a+JO7Ph0ZXgBIcfA3GDpHkPLKIs1NJQEsj8VI9vv4plMkx51vJBXaVuD2LKovn
h6bcBCCea2yFB1EHjwp+n4AR2BjuJum/eMwlw3Qr/1GzQLteyq0I3lNSn68/8r2q
PZ7ocUyqkSztDfBOuUIDtu5J7RuCJJzdpjAdcZ8+4LG/k/M+0dxtUX1PFuTJvO9g
2GLQWR6jlXLt9hiHk9Fiv3a/04qRDVJ7v/+isHHHdiN7EJIKsexIElgTgNIHSENo
pksIgKjDTv9ss9IOTIXl2pgVwvOJ5rcChFHV6cQVkeZQ9+EUV2ta3RTpzwwpk+mT
sCupT+tei0V46VGx6Gd6ECAeFHnOBcoxFO3ITgkkJZnR22N26tGcwj0HuztVt0E3
zjfvokGiFEhs/U1cTS95DvkSWf2KQEzB6CSlaXaNU+tG9aDsglq1m7zYPlMvs0o9
dlag37pNkTZI9eLataMALLV/bh9jVirXAtdUIfP2N/jD5ovX27m23rspbp2UBGUA
uOOS2c0QpQvgjjOWWqS5gDntvDymcvDsDJP2+STCiCHqmJ+6+mm2o1y/NGlgGlKy
NuBTHWF2WfJ60RGRw+iAfSjBHKF8Tr/p2e9GqBPq7bd0kH4e8UlCtCB+Hbervaoi
nn8h6vtbAfqMKENdZNm97DrsNneoRB+vGTxrbsY5w4VAB8iNO4TOWLSHo4oVFx8Z
Ik8baoV0XUVwSflhyhA9xmdO+BQBMAnp8dEqVC0xi25+ncMrhiM37Z4luIZdOiwM
pqP+IKn2U4Y6zPNc4RjTXz1cM/joaxSBd2/tMpjRxFD5N4/enfj9ISW2YZV+uJyV
0n36bcCcIFtHaQZh6XwgmiyZbzDc86xFcuk0xrIK4glo3JYDmPGPXMHOftcggPod
EAs3Z9LAKeGBe+yNlSgiTzzSldb0r/Vwm1UI7+HCdcQjhYT7PZJZMWYYx36VpI1b
4RfjABZbCBhtzhQdFC37qUbUhOHia5YO/4iWJ3wiZfabUyjxkqGBxV8/Wa73ByTI
yc/vQrsSMZa2Kz2RBLRCRYuYTe/rPa1SiggscdtM4MzJffsiXgJMlfL0lKa1LL4z
UU1xMDW+9GHgHGbH7edjoXHNHfpzbdMd+BEl1E5xFv/HFjt00HWnkNstxVf5XuPN
JwACZeh9JpSwOENy0oi6r/GsKZPjRSGgKaCHPSGU1n+3V4AlvIYZRIyef36Us7ok
94GNtLbZeZq0IEgRzRd5HxTbB1yNJPwdwGRslos7yAqQ77vxGKa2Ju2I537ENHoU
8QDgFEVOaUnpb4mWab9s4VxKWUbFWQqDqS2kJofCNfgqp4nTWmsbP2b9SxKh+1zt
Yc0wS17UmrA7XoE7L46FH2NutMWwCZvPhuPkvEBRVRez4aL0WTmEateeFUvxwaV+
1Umz2u9tuAtmeobJBzbo4+CcQ0uyGQluh/mDZN5Y4m1/Ml7XmnVs3y9trjYN5rn1
75rNZ22ZE9UVSX0ValWtL+p+lXvexdCEY7mrbOdMz4sQ9GXDiIdsTH6VhjpXUZMt
Xgapc1173kAE58HryD/ZxQuiv1zWYeCqozcNKJifI52NSaDNodzestDYyjfYhJmN
03Utye8vg/KzRsSCU5fqH1zaNyVQAqKrda1ldupN1HRkEmbZStr2vJ/WrizLqZu3
iZck74bbOrunX1pfo5jIf/VwiwBZwzfPIBpQoDtC6NTxQ6HA0GxYqA9H9KPjALbc
fv8vX80Z8nJBI9z0KYoXKRRbPRkoUBcDR/HwdieRBg2rM5mYLdCfsgDLtoA+a9zC
7zR14/edc3t8RX8z7WaezNrUpy0UPz4hiJrTHDBo6Coa0yCMRWFB+PoT0YgoI59H
Qdj/v1ymXrojJsOfg6axPRVL87oKh6jdAujWRxYF+3v5dqtH30VYxPkY+ERm02+H
YioplesthTOKcNnXvJHJ7kIzktNdOnH1nf2VdZO2bqU2pgWymkOu2dHarfFJeS/j
I4ur2u1Tmjb5wQzVoC6ZqVvGK2Xu+OOcEW7ChY2c62gfHZ9B0myWFfjm6PpNJk1B
lzvYMOqnh50QZV2/2dBj/4xKmTbHKrULO3Ui7AW3LZtJs8nzs2qVlirSM7QRZZX7
7fJ+X5e+3leggQmmHA/l59ycoWbqQrQcGqslYqs3UdHsfq8yMdzX7DyIhQqAFBTn
7mf985/LvUVNoujK2EqWt5Q4N1Gag41L3k2Ke/1Ll6P1PAbU1RoTFEhsI6WAaJR7
JjLPSQGod/Xloqi6QszMkLKKgy7FmO5nXtSAZ/ZwM4bPFL94nx4tVp6at1ApJcnB
GJja0QUzFAH76Vjk2RfSART/H15KHph3ebEyzh1YeLyuYCO41BUUvmV7WFLLaP69
aWL3eGCUGirGeK6ZnmvBMGd4NCmICuYKfBu2nCOEljE4DG5ckF3EMsW76G4ALtZ+
/8xPMFy7v4cBAjHRAYRRKl4OWbN5WLRdACWhMItEGmbAxZWfrR15WnrKxKTbmleZ
uGtlNkaRuqRH823PAR9lB7RpLhUH73k5zh/vwS2vWY+9jZ5wzcOsVI8PWONvUrzh
/7guvRqZjqpuI0bBVlWke/xymjxaz8nWtWX/wmyuaSxEKxHlV6ZsfGjOHtC9qqq9
kqvtphespPh1cO3jHcsOQaaMX8PBda2Mq5juMJS8WzIZIzh095HK/7/6s6jGk86g
LTSywlj2DRJTK9DR1xVMlp5MlwQhSt1YQ3Kdr53HSbuj4B6M/HK5brBBkTG7HyNV
+u3jHARwjIEtOGny0OAPBjPjK1dLwU5pwbkytc0FVUzrG7wsidDXNj5NNe6ZBuOU
8XvIzs3te+GCaLy1uRHK42lEJxltdzrAHHUm2C4UZyVsgRIC7UX4dizWf7b3qUTy
eyblkM8u00fD6r6Smz6S3+u8I1Z2VOIMI36hbsHvyHIrFzcCIMDE8UCY3gqycNvp
3Czx5frri+PnPJUC27jIvHSJDZ26gQX1wXNhqf6TTowvweviwJ/QPvgMLgB5YStQ
In3P2dpTzak4nypGz5VmnBX7887QQQW14ywkD3KTtWKgoHTt+Qe/jkrSYzzx6P/2
hodNmbjcuy8KiyDQYxRwCuXmVVm0eUs4qx1DiQzJMKtQQP7MPv4GJYwp6S7FYLKv
2U5f+mn5dEf9WKCGW9DOEGebRtcCUK6HS8drp515d9gAPw/80AY1Ko4V/Xai8mtb
+SoBUQD4x95mxQxwbaSkq8Cn0ALFnna6oYc9tzDHIEEKcSM9K9uTRBV20mx0ZJ0Z
YAhiwF7DsSK1WFIU2wqF6pYaHwelf97oDNcIeyB7687zS5dM3YbLk+WVCoqi30J+
iPgKViK5qf20KLOlcoRQvLTV3ocsjC993k2KynPJvoZTD63YlyXzrHs1JY1bTgAU
uePv9HB6v1C5TPZcf9UyZiPK1NCh1Fi5lchJQXAMcPKusvAsLcNsvplC/4Owhy7Z
ICtRYL/iATOOvPUHntmiRuYP1OLigbDSFFLbmj5YLAY1G//s10IGW8boWMXms8ZE
pKxkUljS2/v5CydBPIlq6WqxGCHs028eXdnV4xn8E3KoaJPmsmX9IhQCNvtgIEln
XXFPwnzZyHhi+i9lKYgm/BjW/X/k1unOTcvwAPuJgflvR22DUrGmsIuxa12IoPtx
tZxYie9MUmfaHK4GCInvPkAGXoBuffmD4H0KRfM3CMP0FovkSf5aweEuEtf5lr6Y
+DQTEUdQ9HCG04ttqoxikA7Ab0d08X4QsjAHKLO5OmCXRTSPosdR1I9gidSovr31
sYldlsMqqc/d8ryqhVstgMvKTOcLzzzfl4WY5gCAU4vSvTQQ8MWqN+Z/tWpEs/4Q
4qgpzpsLk3rxAJDpbQMrsTC/pOQ7+ZV9dfW8VVCmFUKB4eVBJiEwaSAPbXf5Iknn
Y/Gsl550o9EhtyOwRciyEKzYgboNx+27Z7EW6FEpA5YHfnTT9GDnABipMkaIY3r5
VIb4g8GN5alp5APfby7FY50m2i46tGodxZMyncRHktY5jM/rHR+v3mXFiN9rqhQU
5e9bYz/+/xlBK7IUD0v+aWiIcxVlzWhKB9S8UngZ8ujBOu8y3ci7ALMGgo+wEQfR
4Z2+E4+CQ3O4/3mBzNMAnyAR/IpzqWv5JpBbGIP3v9Lnmy6/mh+cecuTlvRnIz4r
i0UIch+J5Q9QDz3UnQl6HJUB1SulGL7Q5rw+jrjLY+3saOFItacq23WL0c2FbtXM
2dA3ndBANQpSL8SavMEueTXo5MTKBJv/yP0OEANCzTZ2Nq3p5q4ceQy2eWplKcp4
aThbh2KTIrVFu9Agvvd2d8FFv7oaJcdi90RE047UsSY6mY49ezj0rPd6HK9s9PEu
DenmNNHwv6IkzQAtLYwkEh/T8Q7Zy6t2yfOBve/wN5y2k9X/WJ1rYRBkG09I2BKy
7LqeO5CglBvOY+cMW+h67PnjKxm08vKwgqhbiV1aJVp7oCWZCm2W5KdBuPQvrsu5
PkB5M8uVvkbn7S++HSAM9ZvC8u8zvOc7yd10gDxW4EB3Tv2P/+6kqchQ7Ax5qp+x
H9ovvxGTzvZOVokuOP979kmI44FppycXyZyWo9dmA+9Ll8UDmYeW0Nz44KeCGsgl
aXXTSuq7Kf6ksmHkYorqoaxa9hAFnw+KB2m2dwYyhayVx1nQoMnLCOq+oubHgwbJ
gCIgLeb9ibPFVBAsb8WYkB8mxUY9+NNS+N1kKJavaViv97DQ2lZrWWIOb8zgtpYE
4Suv6SQTBAkxz9WrPs5SBwxSk/PXyE7ACtEpsD+58xw=
`pragma protect end_protected
