// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:47 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VdHt++2xIzMMokJyYxL1KX7gVVx41M51rFfKaDhFAOacT3hI1m55toI4G8l1qidR
vOGDTohEjvrI+euI9O/Dlt2TxwG+5lNyRllqHobgCSaVN5xqmdMDAgItSpdkdHIT
DAnEm9H3p28Ic6o1sDzKC8Ssoz2DmGgeM71ycbwGZAc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8784)
aXjSxgKs3oWIBMj4ykAYRTgCCVO9Sw69Cq+tOXJ8vWjfEeYRZUb8mAzklJBWjhtS
MI4GkELhsfLGKNcYdke+TB5OAJJYk742jE2q0Y/a4Kb4ZIYlUG5vNCaqeKK8RpaD
6gim3qwWJDfE6oR8J1LzxGGr3YyyntL0FXK/FQXC2LtRG/eh/4Kqngqcy/pwZF9k
KqclYql634camnQhU7MOZSCgMEp3KdWrJ87Xc2n4JU8uaxFozwJW9bd4ldYXsW+N
g6guZp0G789oq9cVUAioqHrhTm1cCWRPMsiAx9gdI0F4ntJ3q7mCnhb/Pk/7Ps/6
EAqkSGdvikhzTG5wTO+EQc7vvhip7GGlLXy5dDTraNt4A+76wGmqnQURTNILqucB
MfFw7vEVSmOEyeV8MWRxwwDOkC0gRFLnSL2fh+iqAkZZxdorBYH6ZtCLJmYZ9F4M
ItUE3gPeBq8He+/gMbFaNPrD0J9TI+x84dAasEt3bMr2QYNMgE5HouBXe9qzf0KL
Jz9Az+cIwUiLDW8AnIPy9PHl6UvPfmYScu1eIpYstSZB59x6fn1SMJwuPOdcM7E8
sRhPipEe0sYYE1nNZcRpXP93FHxD+E5CODRpudtxHfUZD1noI8jW9XxJmR7SjE/6
GJtumDKQC22fAkQM+QXC2m2elnwRKKt4znvkblacAEMFFQtgeBXLpia7OynJfOPk
+8Bm6QeVQEVqjTqyD1hiWSfensW4YEf5EQWOjqxiWB7YW8vgiGf0zsbYkaFvGx2t
hT8Ox0H19Z5OUDcZ98EmL+6/vSfb3YxkIoOyZdrHEhFC+fRYU22hy+sKtogcoKPW
mAUBcC13/+YEHjBswa9ljJFbAPZitjdaE9d0t75SiPmBqGb7ElqdZYdEvffZMH76
R8simN7solXmZAV7qnjiaYyQ1K5Z57AtncI/tefutYLdro9h36v4cS5ZFjzsGQjn
mX+tGIZYgKakpy5GOn/K5B092jAOb7VeEWs7rs6+Do2pe31HJW0O2FB+GHTxfhbB
BN/bj1dTzekA/W/PpJciQq4lq1EGN0CwoxMhz/2gGycEPirAQl9eikNSnr/0CF5Q
gx+5zAxVaV5mZwbv9xm3S6jBykpLGNjkm1dr/MSBYsac0dZ9uDvVGeqxY/XbpMFt
hyeXudYXztm+8b+ba9X7TI3nBAXDJeQbXRKmD84BBv/bZMMuMTQ5h6vsCIZa8A37
wXnitsQyqrzFiK61at16GUFWBUYop20b9pVGJzLNUKecT4AXPU/OHB3nXlmIwk23
9ZVBy8lh62iG5n1C3cGU7bR1LJBoGhzbHrth7roxVZgigI08edg5QVk05QTg+4dr
M0bw8vXLtfBN9ih/Sy5TJChAWjH0lptKuwfaidhuqRcKuK9KZBo0JtuyBT41QH/9
u+MkVmaIoWMRe1TwdwmwTGMpuk08Zp0D1EKE3RIKSCGHht/sOniVw0gEWnJyKHW5
Jdw1PfTI8y4MOdDvqz+0+PhS+nZ1pMEHbDZZzdszzNNrNs+BgG3XXqcH+xLcBnMV
rqwtciBqCZoUA323ohF4p1nP21bsdg9yR3p5VdtMYRueTiv6GmJ+ovXkTvB+HmF3
7Lp+3BnZJTRWYmrM7fRIVrRW8X+IGO+jLt3rAHdYqYW7j6l3OMsMXpllzHL8iMoN
dRlmlVZrpOq7fa7ASUOpoeJ9jcNIVz8ZyhkwTvwPDT579etPZEOR0HuhCm3E5JUd
k2wQ45XvJpZ8EW1bHr48m2ebXvdf0vNUTYXEB3YwI4k3zlw+JPLz1fgVWhGuC7Ev
TSN8AAkG0RqsSCYIfiZ5Dn98KH7/luwLeDz1ZcoKNz+ttEbuI/4Ugnuqn+Imymzd
CUainAwDVIkc+0c8V/z+RB+djwyshgIr+lIVjuY9hwHhpj9ckqqUy2epwrBsXt/T
lnvlt60Eux09IYO2g5Z+6YA4jAoatcP58ductAVNC7O6x1ONqnn3Wouxs0zefflE
qopej28oh54ZiwwHQNZwUntZrQNYuLhBzVQVppvn+P8zdCnxrJr1olen0l3m4enL
Nejs/+/yHczX+8gpQpfxgrUzDoZ2Pq4sdPdaMAFN+7Lat6EAiwOcl5L2q9xlWLq3
Lsic/OOhVqIhIqAfK5HeBzOEecwzsoRD1DMhjr9MQDxXbKtZiPvI9yeYoRuSSvN1
kRXEO62/sypjFilqWCgKznBkpniBq5YG+iMOZxRzEBuqWXOqPqVe6jZ4kKmRRnt6
quQbQD4XY0+pICS9vwPuglaaLZV3efkNu9UNz8z+TuAi2ZJqAePSYQMyloWohc73
Q5UvkjaP9OSPmE8DVkXv1Ex4qRpLnuQo6czTuZKLqlBAo95+SjYGH6daKE5pulVa
Ny8ISHcEz73Zet2PrAKdZ4CU+Ya3lSYPQoUebJ/TUtYWJtX6zzotOYW/PwBMDupd
qXaBcuKRl8pZkddZUrso3kImHOAAFHEwe+DptIRN6EHe6GqfRyV6DdFiLLFm1WOR
HS53ajp6L0LXErIudJ9LWQ/2SzwFjbOOZ9QdyFDJ3zXvh5Dzn4WBbtUCNqLxY8gT
O5EmF63q5fw50syG4UwNm8j4HVwwW0wbk1UQ1ao+SLbNW7oc32a0Oz4RkJuyVb15
MDnUIYK4aLf3TZYfVQiMMMYlW1efH4tcY0Pl1H4SotsW6BYnaPYBUkk5tieXVia5
+uAIp9A09Kttb8t7+CXiRREmd64OhBkom1RRXVvBnuld74Qvx6d2ChpEFNjBSkg6
hir4NIAvlJZeBN/5KOh5nK63bYgeyRtwqfk5kH1QPOg8fYkM/Y8xipTvPOYZFXi6
iec6Bqc+tbg5yOH4L5gPaoy0m7jnOXc/Un5KEWUpkgHSVagqmn4ho+FIh7Yh1umB
x674DovumPbbaMPEmunzqt41qDkwFQoIHu73kQk38VAYlQtcFbr95Ip5Q/Lcvrqr
CSsvxUITKEjEF6wj90y9L7HVtWokBGSdnhwGcdubwPj2mV6DFLJWfyGLkgcq1o2L
fZI0mllqYAl1d8bgPDsayCcQpxeVDErGxFc/C/6stoEV0klvFeOFgOcGWrcVC/V9
VCriWG2TbCP7CF0Kh/6tg1Z9npppVoGvmfRTNs3D5YjOtr4mggmqPl0DH9DKMjAg
57sao5rWRCK1ytPoLOkJK/qVHlj5rR9ZxGX4mVziBhKQg/GN+txI13nVSkDwmA1e
V3VC1qrazEyY5Jp664IC+rzOrjs6k+ZtfdWFyjYJkM6sSWGmqUY65452/PSoEehY
Afe04PD8gZuCGl/Gf8c3JynAy5qIoE0haHqgpiBIoYGIkc5F9+CWH75ZsJm37TOG
gvpT7r+iBA4rdtUR+mhxnbSpkKz7dffJy0iBmBgafKm/+nsOJaR+JDVTJPNH0PLH
PjObjiOsEm9WozCrEgQFAEcert698Bqk/V7Gq+UMP8lSgZV890Obqf41h6oaXNTs
Wl2FYAsqCayc1+YcmWQs98Zb+8K57VBgFNwKZtI29OS8JHuZRuCVbSARJuz0Q1xs
z1A4GGXxsrAGta9X/0FtfVe4zODmPr5N2gTH+A1peVL+B9hXliHSU6ApfJHab+f1
4jEkbUNO4w5F2LJ7Z70N2t75i1QiN51XcGdcxpyZWfxoMlplS92SdKwfgOJezzRN
WadeM4xo8fT2IWaRbXU5kBrdEWpBNnV/u6o5tEjlHNJsKOZGzRoXWFKxSo3gtUr0
ySMgroJMUEan8LHNOymp4oaWd8gnDGPGnZsRhLhkcpBoONjuA2Vk31OA+3N8UhU4
+Q/as+A7Qsi8aVaoTiDSJS6eQI76IrvMXvrABMJuhjwpauZmUm7JNkulFZvSi35i
V8s31fRURmfWp/JJ5fsGTFEhwzG5GegkYRO1g682b5PlMAvfRZcmF1VIgLnfqAPR
HUoufZ2OSwsgpG7IF63sRdykhdUY5RV+7tmeJEk3EL3sxeAc6xWEjOUDv+VEczor
UPiWSVS8YD8FxCtH7Q13YVwCsOdTeoj+bczjE/Z3ZeExyuJjHLSNWWCFfKG6eJ5A
nVRgm67jMp2W80SkChoe8mfbpEnKpG+fcqGNDsOMFDeM44c/D2IuPDpfog2WHMO6
FpGGRSSpobRcn10Gyo7MvObquMtXLXhDjvaavo79lN0iDgIlhixQVAkJr4k0onr5
eOnkZXqW41gs4ZujN/quj+GX8DBcxRNjcvawOWd5hs2P3I86cRUjr6FhU9/cZHzH
I38GFCvgl0cmmNtzuB40kf1eWqO66giPpzTyU0xOv/T9CgawXch4trycDXJBK7x1
tW4KasVYrE8Wj6zlimqDUu1LG1ldNCU/lyGbyjlshreMHnc9A9a9W7w2+g1LM8uz
VwFwSl5qV365c2V5stCx1MRFz9nfA8g0Py/ZEcnHtvwUg1zOgE/Tx9R5RBd50IIb
TfA91srsXgtCrRbgK31FKsZorZSls9E1MQj675yvoiGDrw5WLanVjNGIuz8Iccdr
a6YVOmLvLjDYpvgizx0vwiOw0Ve6htmpXUMuOXihbTprMCHpKKsu++RedWaQCdo0
Iix5btsn4KLHfzmTCLcSubmn+NSKZCIpbYW4u860h9cDaDDfa63lrTx+T3DPCDR8
ZEw/Bk0R3wxM0FbVnmeq6MOVO1zSnTtPCK3XxMGUktJDITJvSrVapnz6+bbuUPZE
k8MyGgAAYdytHXC6le84cHSfAjDuHga32ZUUY3KTEIl2lkQNA4ahrIx5OaO0AUpn
yzxRazqZ/gqtd95cYN/YdH/oSwokpQlW/dkZw9y7Dh88sbmCapv7ABlBNKE7UdcH
Y7v5V8GYoEbd/CGbbWLfTJlRQdUk0F9JLMrJQkZ6RFGXCPpxM+SjjYGJ5Mn5QOv8
0KvSzuolir1xZxrTaUGxKQPMFGgYAjZBjfLnZqcxeHIW8wM3EByeOd2an3lkxc2d
Il2vPW52oE30k8mZtN7v8jLz9++smMT9NoI5TA8B2zFWrFNw8TyKauTZec+EhxZZ
v7A7j0rqNsegITOAzTXclJO9h4j3erLxK9amAOqMdP/moU+qfaINKQBW8RTptlkv
EV6MZ/fMrMmwLoanH2+wWf06by+UKB4uQQ+KSDU8O16SNIT4zyEEYYTK/gjn64i8
p3cJ8LlzyIK9kkgG2E3JEYgIr/97fimGN/Yg+9jQ3m4/4f7f4wwUHkcFSdV76ARy
BgzCkvPeIlTaf7eSqfQRoLLmWLPoTABlIQSO2O1IKENi97NUFFUdHtmFwSOVeZ2Y
VYVmKk6YYkGy3d3ZTY5yg6W7ogq9wl+cVnW7vuelNGfA48hcsLIGhEQCxp+fiT4I
hrNuhYkKIxIW/A5TKFJIwQME5qYDeeSu0Og8f6HfkZSNb3LOpePdIFqTDu3qmOFp
BXHeJAU3INUfZUSv9hlC6Ma1F8rQgjqElqPHQf4STtAysQIBBy3IoqW0Vgui99OH
vR2+3C1izPQyfE0JAXjdGfSEN4tBBA9EbQeSCaPy+yPRkIptj7j9pt/GamAgJiT7
zLpMwW6yLFcYgaekSNuP2gxO+NsgIWHRAPwmgBbrM/A4TLTmn8fQI1Nl+82vqoWy
F+srTFRs770Iiv9dmoR6Cn91vXvqrrGJmSzlkRK7v4kpToWI9ZJ3B6xly2ytPVzb
IFrhm3n2nh61ZqKFXxyyGcQXD9XaECQ8NfvM3rHWTzg5vn3U2KzVRAS1/KvdpVIe
EGQcVki12HoIZNk/F/KQKDaXglm6E1kzWMklHjBh27RrBwzK3U1QKy23ESO5OfNU
NWfF6I2okAmksBIoDK+kAyVfPHXXUE7NqcTv5MY45xErb7GL2yNfS4V+bjFLVOHu
LsKtQ2lQga0+cv60masjp7zesjuKaWEjDljbDK5tH91E3acWwVdKW5serij6YwpB
3tADPU5M4SOBnQ5bqMpsJB61qIltbkhOvZTJFap1SWOBF98/xLmKN2TEYWvcewD0
Imn5fIGRl07pAPJO777rDCazd0hSuwyVpioxBjd7p5P7e/wPOdmQNSUPa5ySeIzb
YCwhYvu0uc0rZcZEmgjsPEUqDldnDTz4qY9pjqiVSE6xK378dqSJdooeh9RwxMt6
P3lU5cDZOD8pnBM9LtAlDf13zolKtFnIJsb/IOx+MGPgWVDT49MEYdvqSXA713em
KjUnTKIRhAX0OZecE2oifHA04TNb9jygzQrBSF6eFYE5yT4sDTYWBxN8yn7P8U1+
id8f/dcOehE+E4dymIRe3kxbgsYLbs2mWPKKUBTxa102VXHMNqUR0uiStAnC0zdn
c6GMmaNgmKIciH//jq1VzEqmxSx+kvDA46oDCr0QWXB0014UpirqW1l+2T8UhrWD
eQ8zrus7Fjk6j1+jHXJ9ARKk1q8CljmuGA/TZaZ+XfJn9GjbnzoRrxKaZsZHpyte
eACER+UJDG/RCnnbRVZAEGwtPJrMvLh55+2ncYIGBlBNoG9+xLBOs6Ogk9py+2nI
F147JuV6e49Tt6x0t4y3fEYUxZKGUuVXEZ7p3Ljz/f1k7YtPmFK0DFDVx0vkX1XP
On4htYF2E6gzUDM+CKs5vBM9KCiRr7XulMvWVzLFoOr7tsdbStCheOneMOTyJT8o
F0F1FpSu8JK6euSXWx7iHpgTx3oExfw0P0pt0hK+EgtEJE1VFvhgtb7YNBTJPLpw
s+M8NOTeJKLUNT9bitGrmDVlz8VzC+gC1MSBUkg4L5shTzYOR8elwziY9Vks+45l
ihAQXnNC4y2Bt4t2kzIZIKUhSwZ+iTr3NsWcEe71UELcq3Vf719xswLVb5HRE/bo
DtoXTYgjxWNZsBAnAwPDT88kyYC/CpAgBBSu1Au2V9tq3iLouqGewn6nm7Wq5gBL
drDQNfa46kK5m+pAwtvXAuMSAQ2HpTjp8Vux3aWm09hzoxtxpRLuS2ucM2AiNrpu
ql3eZ3juqq6SBzBe3ijoDGu5LRcMEmnJge+wksjdC4DhVeqMixp7PflGbYn36Qte
bTvxVJCoFw01dq/Ht8XQI8Q75PdB7dJQ4CzWE1xm4JP9UYARF0ltN6t27VQy5vaK
jYVfzVCw08SAV2oJQEeIPVoHInjNZZaAcZnloO192AmIHZoTRqZAMSU68TgOQOmV
gsG6EeuizhyYPYZ5rD6wdePeRDDxc1I5kARt93H/uFsLyrdAtV412/ToxWW4BDeC
BNoI+xwiRlRmRxzsDN9GUmCHm4Q27PAjwWVSH8NdWkh3rmTtc0PN6dtxSgPth1dq
YFIor0vZToLYNBtbblf8ret6loHUvywBoJ5SqwoTx9+nMKksmGl401rkpoFBOIc+
d+x7A9FbosjcZ6RXw4ZBPwiaKi18qZRjVIqTce/oSq51ghtiEE3xKj1eeaj3+y9b
2grf7Oqeag+6gtSZKGyMYv3hfZ1vqbwMVBVKzHm/RsSIZpRv50LzjFYadscssRnh
KVYDqGaJyxAnrCotWObb4zG9U6MdwXsoeByRX5YFfIBL6ROWVXIpVxzyWahEDdg6
kIGTkBdauTXGyZ1P9hiBkIy4zoyTZv6OOEAl51sLmGk9d4QxUV5wprLoTVmc4D+W
h5OC7RSeL6ZpnU0XSOfB05bQEQgMU2MQimCKoBSMLToFSmqmfDMpI9K7rn+Y5G9N
8QhakHVi0z8gkwxhMH46Be+QEXVBL9LYR5iG4S+tbgWbxC0M9e6S2UOJkVrxuT0c
/9v1qTD+5+LfPntCt+opH4Ekjth2I8QkuPpXgsuNCZF0cqGAYTjsaMRJzY9gclNg
cqtzrAShnWs7EyN9D3v9Zrm88PlymLUNb2E2jpp5TfYEW14gqj/tOkWwGJlctDmo
VDQpUopTnf49zwnlKpqa9AuQfKNChUQe3WgtPKLR1VaM2qIR4b6v6fAfevZKRBra
ppDy8OskfM2UkRNRFreus03M7CJTUZpAXy619K9s65QAsi16xIfh/uD2rEqv8is+
XEtjSLmFOKgjHdsRfq2SKwV1QmcQdW9UabszGY1GHDl9fQUJmgwctwvO2oOyveTs
9j9vLhqRUFQEmv5nNh5yTmWY5THatzAtO1TSuzcoaLiHsIX0omovPJMkBjs5IRCN
aA+YbiOFeIAzA6qC4cprnmBVN/PKrUCoE2PFmI5QJwCCaaoUOc4mCUliMRWxjSof
t8sU65FAtsUH2763L1cul7VQTonnzSFuz77222Z3pFncIGODiwF3UyGPr4GhzgjX
nQP05rlgcw7CkftWcYtl2WjZukWZGI0RkQwsd+kcWbLZHOeYj4wRaMfXmgRk52nx
P35g0Cf8kzowkJv/3WQWFMcZYcOes4BXAxp56ipY1HqZYCeqKIGpvb5PHdnjaqoP
aIABEnYdI111oxHmTEAQZI3IYyp+9OP/1KNKdx8dZWa/1ch23hBDD8BBO1XgN39w
AD8ee3I9Pr88ey1mvDi6A79zgYSW9XXBxogrdU2c4TdZ7Wzh1mruCqb5hyiy87GE
XjiHJCR1Yeb6+KYeJzazct0XsKXO7lLcstMMgdw2jrHbdC/ByPimAwLCjrAPchdt
ZRGnZ71SboTT3OIVtQsjIXDt+eBlLFl8dueWFpoadx/M7omoaX/gLjrfMh5NqoUp
DhDQKlzytLMnW6zHWuxV2Y2yAH6Xe/GQij/1NIgN1HsYBcv01wDtZ+rPuFFkDc5H
RjfmCo3uhOfoiwzdNpCK8ohljuTFXhsvm+rfWhheERiwhsMQudHqNWhGqi0wYrsQ
3YfYVAQehhBmAeR+01wloiE+NdHkJRuRdyvw5vYqT3OKIq98aR/C9EjBoGqUu5Oj
AN2put6tvc8MYSTgO+EPm5V50P/g1DEgQWk86SZwzGS4Ruzv9HX7cDY4ClimcSnV
09JflNv4n0PHkXOTSDY69cdgMmBKve4wS75o4nXzW+IVFETVlrXuZ9JXbUw15Ov6
zaaq+SuD0Pl9Pc7ZPbcgr1UwlxbDYbczwRy0dff1VSU+C2iUkO4Ce0w6XjDRekon
jrZtt+PKMeULh3JG6Bk38sHqkf+m7jzUm/N5hazUaP6XLIfkHQQsrdgvloGTQHG0
Icwbp2ZBto+pcl8KTeAbxAEzlokiN5huZm/KSvSbOoGBfsXvdiiCqDU0AKkSweCc
af+en2slrr9m8c73kjgbvdg+FeRmwqQ6N4VNru+0xsfmSJYDU1b/Lc3RcByxi7Om
zzLrQZCQXrmSxL17ceubNKY2srLCAUXYB8JrPglx6I/FM8qiheUPEV3yWbVZ9VuJ
g5Owl3rI7CBkiIBPAILAL5FJhRa7r9327rfgF6Nbkbhtr2gXKm2wCZNGSzz72j6j
mX+B6YOo5ZjcRihcIxQdN/iXty9QV8NTx9hEq/qUrtZbaz0oNek+b1A5u+3TU3MS
xNHqPEiNf18QHawR42rbrQYl6Zs+uy0Wz8vnQBwvdsNDl6EOUSCoEzcqNb3LhsjM
nWIKFS8dzgXowgAn4zVqX9R0rcpH4wlf50p6WVmtQyp/nsdTHwADbp30Bv21Sads
b+0GkZzGHC1V8pYkgJ39lDJfwufWvbroqiYD0u+vWqFYMmPJJ1EVKtKa4b0DKBlg
USP7K5GLFyDbhoiSSyMDDB060Q6kYvRSMi8AJiwT3JLwQoftTfEF07j56My/JGX5
DqW6vxMB5pIeSZBEEyBlnF+UcMt1vNPN7ud6LKk2Jehp98YFBnsFQnp2cbZM2SCh
6BVbSKJJY9ZeGQoXbNGNevBv5crX7EJQ5QBCACcluuJmWTCRZZ81DngxWSdZfU+5
NLOKvvT6+d5CvGELHMqAnhEM5LF8oAyyTAn7aQs9fHb9WkVvFi6gsv2VX+yQ/1d0
AHCdyKPl0aAIyZ7praUdSCoUtwF0L3ISDY3S/D3+GBIxblRM2H+S+VFbnecqA5HW
IiMljxiReKWmfniQhsfVl7j7ni+4+6sJxTCJUOli5zGzqVgzayRkv8MNq13lLNdk
TnCU48dUw4w+WpqhDV1HHh/anPm3EBulXtE+ydfcgD0BejvD2QO7HzqQBPeJ8ZfH
8IsJeD1wSpOiHchDvpW3FF4y7FkyeUKo58O1zC3AqSgcnvGzlnCeD5Eqc3ZnV3W6
eQWReqnud3r8lbnO8TLORx97uHzrjqS6J/kXQEcNLjyBE1V0Pun+e4ybQi6xidbk
m2neGfzuy8G/6IWU4w3djX/ycyV5fIt9/dMlv+9UUDOH07f62SAmRv9QHf0yFuiD
zcYFU4WGONZkTj1ZO/4MLDyQvAgz5S2OzVS4YQkqA8FlwdEV3c27Dvi2PRu4MY9i
EDK+QUVG9pqoIf7qMXNO8jec5KFgUSmJrmyJJlnfWS/mrig4tUQiTe7f+lT5AkLr
IuGl/ULPNXxWMHK1LWy3T+X2ccAmQYf1zIKwIeyuk4NHkVoAfhlrWlXiks7MEHhy
Z07SXIXMWSsmaIs7edT+fDofORgRjNNeDwyxbbp/jpDtNdn+0xrvNMH/htS4aTX6
ZvRpQuJgw0xTMxaBvNrLMMbS/lqQ3IH1EGzSw2UYM5wmJIv9ikC+SBk5HQm+eXHH
/E2lCw3zIShovudeInS3X17f6rSdsxS+Nad++WBCEgXEZstx68i1MHhgkZb68qvb
2Bl2sdqiNwT8vQlm9jNJfL+wpR1s/pPt8TnDOJwzpbiLwc5rlegQHUmJsUtSaUWu
fstQqYc6BflSeZ3IFrwqorG3REhTDRVh28pnHiMstUEI8G5Ck1S2ZWgc6QL8U77P
5jbEzYtvkIqGDYQ7GoDWdVbtTibHnEs9soFcxUpIN5FvdhPX927U1l20k49bqpkH
hePOWy4l7s4RM1gGUBNVQ3rzIGi1fp9pHx5WpefAhJKzLw5TDTyseULjyF0csnpk
vs/CCb5yXGJK+MVcWcTCpMpi0/6tFbGbW7kCSOSyCOEo7avyIogg9krKapt5RJcy
NLxpibyfghRS0vPdPEs+1hKkUro2YJLrFPsPsh3ICZfmwVR4A9VBpMM4QwgEUcjM
7o46dkQj2Iy/Xpkf9JXZsaUzg6R4hfi3fwRHh9r8QOxgb6lTVipWQ+kWbJFQDSbX
TmXsxXvVB5pJeTjBnB3kIRwDMCMa3fvshMraJhdMKJeHCmBAN7MqDVti9qKFhl9r
jP/BOLFcptsb6gj0hps2aTTricnxVy/t3Twsa9UPuMaoQO34wwk+2oAhfQNc1bPT
MC49JcESHXTCc1RGP9r00w+2eQjLQc4zdBizBNyypQDI6D04jmZjSZTQGQto9SNI
4iWRUq4MYIj/gazh2nQKc2wC1AggOfIQZ2+GYlHhQPpkCUCnvsGn6XaQVIzT9dcg
oahj22DT51X93GVIrEf38NYQBgKIbdxQ34WUxQS8VxrNSP697zphKM9YwGDyHhow
fUgxKR4B4NrKz0QPUfEtW9IYrBYYGBzVzIzP0sYoCvOoWN+7hZ/TyhCbFHfGJ9na
ILkPgxjs0nkqF1R9BlVYXJ48iLEQkZwdrjy+SwKasj4H07GUJ6jVX6AZKLF6XJlk
jUBdlRXlHtaQn0dBEQV5Q8+PtrO8HWBt6xIt1tClbUea92X63c7oAAeexpSLwqCh
COY+ytqgksNnnrXAM6em/8AxQBYYZlTcHT82l4SXqEPjxsD2nj5gmz+PzzScXZaM
xCLQlzekio+zUljngYxHa3vjtKDeBdzjOcSfz6HB3sjwslH0nLd/h7z0WyKiPDWo
9AqSdAPhbNywHY+lrAnAPuK0qvDw+Hcqc3Qdc1jiKTTDS/D2lZoc5Qe4xeHj/TnR
`pragma protect end_protected
