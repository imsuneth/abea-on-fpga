// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:59 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EV0+WWGNHJgCrdJozNHIZMtKFKU6RekZH3JGF1135ggq0hpJAhpX7h6bRD3Q8rVr
p46MU+qeDnrr25sjqtkdVJOP5UkzZ/9JTS+RI6sehynwxuQ1+sraLDlCljL2C50I
UblY/q3EMgGfWrDORg0Xzs3daeJUxGGjhqO9ppvCBWg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21744)
gx+8SLn+mj++9As88Ml2mKTUBepxR1w7x682auM+16oxgu8jHjmhdAlfrhTZMSkX
P33Oujz21kJ94383OHugPXsqmlmuyY6lqWyXmyOJJgMHWjSDR14rtMZzNt2Wa22S
pB3t3H1tShkPXf6xbzNTRYMCroXA1fKIexIsi4qN/AQehk7CVkgVm1pHusmZPF+J
g12L6EZZsK0fE4td+6D1ewh3pMxBmjbV+NpUBkA10xZ+ujyjDibd39pFoCdDKldY
aoS36T5/cxOzzjzTxvFlA5ZZA6avJ7k9SsItTDiR+9eFU/cl+Ue8jVZVsSPZFvjh
Yjuiwg41/VCRV3Hwuk3LmL+iuu0YNelhOxE7F11cq/xXDe8yIO9ESI6LmSzTiZ8G
RadoK0y1kaR2Lj8GgbJuO/ynL7Qgufi82hRTW605ENxhFxY6p5jZvlldvJj6oOoB
L3E8sL3i01n0ixFblRsRYI2rad921RbF4QQhF6tHO+DVnlMyAh9c23pF0mKw+7mq
bvjnD47hMMP3Boyo/x/AUfa/4bpw13mrLOTer9JyV5D0nU98w2iANaYj5MEEL43r
mXvDnZgQgohfMM1jUnEm3igyOJ08EFmgUrRF73LcFtt8Ok9Cyq6/1i4yqr5y8aSO
8mp8sM9QVCUbqH1XeSsyb6/MOXIIRChh1b1Yq/sQwJqHiCmShVOy1bl6wVG+2u13
dJ/bV/Y5rX8bxtrtVJZAXySHtDC3aw5GKFiYV+8xSo9xV1LBV7PaGJye8AMNM6T6
8KxlErmcF5j0FhUdVNuHxN4rDhLaQWnIix2m+TkS0an0aCa+NxATedaYho572htz
SKonoSoHdTOy8lcv7d/ip9YUlfVPxrkCjDoGtVYv3z7dTjvUDA1mMisbSThnXe5L
/qyXDdujQtbixarV8cfWGV/abO0FgZI8IZdGOPc0L4WbfFdAc2nZV1rofc3+N5UK
JmkRMDRVLA+pEzJyJcbhm6HzD8XHN7qWL4BaQ8B/MMBp9aFWff+gvqA/NWutk1qL
+CMpwFSy6r7pWqzR42z4e231pD7NZt7laOwyXOD4q0mfEeXhSG0fyU4xcQX3oqH+
mCGVXJnnNbvko8BP2dSJhDhLokO8vHe7JzenmfA7jg6Xg2FmlOS9MjjT1omFHOEb
8YAvD642Ajv4P+FOeJ9Wg7shUFXXQQxuFMa25BT4hAc7h2YDv/jVrM5oYHrnOvy0
ZARO/RDjhbn2auA5mVuDYhxVmSrYXg0ai/OrSl5bbJz1E0Xhxy7y5FQdUmf/lHcw
EPalelAIFpB/42m82ZMueF8z300AbPJqGyC2B1gZQFxfvETctDmHxEn8v+EAe2g8
pGWBKg/pjzYi+ga5sJGJAW1OSkAZN8HUMb37cI7z/JrgUvTQ++OUcao9g07nuuYn
Q/z+alZV2NhTnNzwWy3DznkLePYa6BxzZIMEuWhEiyK/vbBps7hqoAp2yg1XM6V5
Xc2lWIwKVB6el3jNi9aGOpHE3SJifHt/l7WgIflthy6BKWPd5cTElOADIEg6yFQO
f1MM6A5JAYDrWAqwqHljrZXvsqFd5fjyzHkgytVzD9wL3o1UNSFG702FMPbrIuaH
E4lXLDMZfEoHJom8813j5jIGwSnUSwWGOe2uNqf0k2PPnLfjg4jQjCPx3m6fBrGl
Vxst675q0Jvqz1LmrRyN9Oo80AkabBP/7VJC8XpFoqVwy2euEjVbKXgws2HWOz6t
C8Pk6YaqWJ2c6jmSbsFSlWJE2vPXweDJ33g0Omip9ATGArRFcqxkITP/kV8drMsI
EOfw2fqlhsusVZprMBmk0g3f1j+Ho6eic3wcjRdf9F+EuDkzn7njXvW9cPz6ab78
OQ+EBrbV6q8GXvCYR9dHu+c55Ym14hv3jcTyHIhsXyX7xEvSId9WoUDzlH3L4HR6
uc4nS35xeg1utq843bRsaOmwbaO7Gst/yowo000REWVQTPs/R+Wbnmu7xFFcG7r3
pDahTNT5W874xPvd4047WZH/YTuZZUeP/Pz9CCP0hSxqXE635De8ua9EZV0IRL9C
1cMjWoGdqFPPoVYiXXAFbHh6kOOQ5XDDPrqFBE2l3j+SLHsdlsywl6TsZpEJbDy0
cW+8avk+ZIIsXs4TpVnT0kN3K4e1md2dk7wLCxqe2mBTjEPP7uN44ms9Dodxs1Lt
THi/rCOb/xOEC9Pv4iMPBHlfZOO080phwUeeFqMdNqdL8W1ZtkYjg/0J/3WNnmub
ebg5IFoV1TWJ3/DIIfD4BdPdn8h1GPjim/akLqZhLDAyZlg/rwdpdjGLSZkuL4+A
DWcG52CrNicbPdLqeSeJVgZmOuCry1HDFaikZsFkyKRPp+85c0GSZclgUyb4UHCy
WDhHvbLuZX8uo4qLLy94rbVj6guLfwgoU0bgdOd7MHdpxiPUzSlac3GL0lOoEnop
o0UmcPiFbG5+7vFut0o3eqsdvyvSozKCPwg3CvFdk2xmVc69mTPSgicZq9IJMPGf
CjUse1lPdm51q9aeujbsOKDXwx+jK67CUahYMbwWYoLeyA2Pk9iXs9gEXTaQ+X5B
GYnOsbJP0s+bhKty11ukb0x8ZOWXGuurr4WocmipTfVFCHEZxyfgZpyYSN4zARot
/5ictCbUqIgF6ufxfRszbRN1pLuZseymMTyaemYYwmODwpErctkpgp1IPxL4CEL5
X11Smf1xeSdOtFgJ4+K77cd9XJmi26v328P0ptKv3haMOiaxkPfULtqiY3OSAdNs
g/l08FaaRSYB34+QD1rrPV+lHe4LQKD8vsVHfDR4QdOwoOdKRZaHf/xylInPW9xW
blk7/hCijfZP/e8e3qoUQWVchcgQuxzvyM/+Fzbqk4dpef/QpGugevoch8KhYBJQ
7WMMv8TrlmPqcGcBUd7w5k3jwxTe0aDiXkRgbWp70Nl6K3PyQ2wgQZgojqJ/CnB4
JjbbE2RaV9hT5eEZsYSr79Ul7WTrjUn032zULaQSY2YT6ULKR2+uCMHJFZ0l/Mxd
vk4SdRW8n6qoLoiU+9nNGC1A1UQQgpiEQLiGU75O8XvFhNqEkCWPc50HazOrQFib
1aZJwazK/FVwK1iaqKN6VvrVffUENQA13E45Yz8+lg2wMUDQ00UMZCwG4OXeRjHd
877rzPxLo35mBLdovQUrX9ZsrGv1yLWjhZoYLBbUORMMzFIu2aeP3LAJpXy1ZSEn
9QAU2W+zjWXwPTjMjeM1/YibFvNqr+H6zyZIEjkK/lxn3MuUm3n/fFgSEZTrTLYs
8S9/36uHIOMhH7KJb7iJfY6tmDXv22PNJNg2en2AtjL9N/Fxen0ymLMFc0ylKy0t
Kqtug6dnzqo886I1qCj++iJliEuWinW09cTfZLGL1ISXTf3E0TS/dcceDTN4jGJ1
xM/2x3z1xKqlqJ2c4DYWWK1KpUVjf48fxBAN+0C3G0z++g325WMnuGtNye3C2uB7
oLgaU2ptpz7Ic8ACA28uHL516Vdc+yZ+Ok0yxAEvZfi2r4ir57tq/Ldjw1aUwj5k
xvzuIShiecTbi5dLryD7G5eRk2+8gwZPG4Fv5r+Og7Wk9HEIo9qs82oDzgMAHKq0
ju6CFzSaVwjTwQ6vPFKTYMtILLSXLt2ryTGSqRJB9zTOH4ePmnMmkmA4A7ppnZbj
SZPCNAk6jDG8o/zJitvved1aJmuMCPgL5uJEoxSoNMAaGYzgYy5PQD2HL5njYzK3
YLt8b2bAOQigZ2MHGXbWf0WyJ8+NRMZ2iFiCSChvrfFaNnOrq+vpMtW3lEMERCSY
vOA++m7LSx9l+tq05UxzDUqFrsBdz0MynDntF2ZjYqkPEPQU4mXxk7yiTlaTdfic
lnL7lQQm7U+6Knz2sLlKEgwBnZNO1w/bSVlod/hY8KiZvnshEAp39d0zr+cykOtI
KEiHmDwXnPrLKGp4qEnF6tgHlkHq4RDmRUmJOJX0sMiFZ1u9VyfzmDeS7aPzBya8
5XP5KTluxW84IxoavGDGoTGB2dM8/rdpKpBQl5ai5th4YZZ4VDObmmRYazAlGlYY
sKc8GSBg3ACo21HRhhLynwb0uj5uNvS6MujvjyPD4vr8tR0v2tmZVTI8rrtZISlR
pWHR6rWoNfu5gEXYgsj6rS3ChsYlBnTIOLGANPDI4egio37WZM49h5ctg1S+fvBs
VdWYFmvmqYi0b7K4V5FR5joXbsNE8HypOjLvR+3lmLPYnRcQFVtzwzRvNrbxvQsD
0OvVobee70/k62pzQwptc2Jbo+CVPrFcPPJ+zbkb4iuqqWzqUQmPJ3oDVD2KRax3
pZSIfW9G+exE4AZ6SWP+410Jo4PoR0g167TSi8KcO5U8IU0Lzlq9s58tgjU9Ow7b
sBmIKCzijH527TPi/LsJCeI8d47RJ5poQhvz3gz2beS76QxOjO0j7yjj/ImN6dhf
HJG9ES9vQaOzQjfm/lpnXd37ajgJz24EMwTeh3L3qBos3tbzTzV4uT+rsLmGTsPf
vE8ZB8CmTjq+4vMj1mB9NhoohGk7CR0IWShgBv1T7eGgrpSGM5sLMVW+Sg87MttR
2Oj6HcZQbJ77z4NnlsNXfJzqgBQ/Ta0gr+kke3sJ41GftgHNA+60WlqQ2rBdLUON
3ns5Pv7LpNJMpyCxg+3NYHMPLnnOtKgs8oQ1xH9ARkCV/4+csYYBEZM9fWW0iOUq
j/qPmlETOTJDfVL1yJvcMcBaodwFMNOv5V5nNVVJjQNqwXW0C0kctJogYDLChHSU
oST1SmjTGONdAJ1YQkxOFQFcQhun/w+9+9urOicB58NEdCFI4JbmrxoqwOm//E2r
qTflJ1re0TIXQmrcgB8lvG5kAhvugZDRPFKb2hC6300lalEBFMSdq9pTAggsQx7f
m2uEUx+nqi2aF2YBFyEKfMPG4n66lxWUCNQQxK3/FysWSmEEq/f9+Q4JcF97yE2a
ySY0eycrQRJ15gCQjm2qVVeuYkvuud4hwU+XQJyd3mCy8bvgxDmEkCwosrRqGEra
MT8+Fovcs0iPPovQbPUpXsWYVGHtakgXMMQ/+XarZHOYk1XIQC887OK00n/+z2rG
hSRDJADnXwLrreyRAGFJFUq/Hv/UGJZDymPkyM0ZJD//NSXwfRpflVKJWbDWhqe3
I9Rg9Z6A9zXzvdM4fCsRMaBjusGYSL4DKVEKuGKhqFdJtjS24BBe/Kwowc9XjdBk
D7ZrKOOvevKItJlSidZgiIaigynY01hFKGNOg//ixh+LbJ7S6q9S/5LzQ+XaucN1
bA9llhiS3Zhf7BWJh0x97cCzYB8n6eEXPkENb/LbMdNo8vsnMpa5zJrMCAHVqIPt
uHqNMho04cSS32o3kOpK9ayAOIPeRBZKqoR+8LbfxFOYUOSsuh+D93AoqcTZuuaG
Z6h0Bo5r3YhLlMyODcOl4PvnEs6C8iIxe7XQSpmEaHAIdclDYgGSFwoBYdQCrLSH
zJCqhxM5II5foTTDarXN+3/RiZx6y+9SCdm4/vr/DhBUS0jJIyFYfD/NwKhVj7yO
qKtsN8taNrrzWi5xscpbof4QQI6uDPKeIEyRk94NgFNQlMjQyMtaHD9o5I8m0FnF
Ff22d/yCFLF5nHR6mQp8tFUv/hyHkmE7Vo3T0KBOCLOUqSEzBTNRL5MgoXF3cx+D
h0Ty4l48vpuKcMZaWMMSf4/h3xHp3tXzuIUf5PU/vG06nBDiOqqw176PpvONHjpp
qNQXHkvgtJEv5InRBHPkhTozsNtWRr2VyS55cPfhYIhAw35wSs2/3JF124ZlC2j4
LVJe/gERLkAPVth9VxXIpFL1iNrxEZjyw/caCsEMU623YiCXLz8vMYK+FAdOs4AV
R4NPQX/DfaJKR1hHFgoxhQ6/W65G0eeHMsKw1aYcz7UaNrhxmdyXdxX123Sp5HSm
Kr4oa7QmwlKpr2W7kU2OlQYuxCp7AU/NqCdCmQB3NLYN1T64tVaucQEKC0PwB6Fl
yC/Vw3v06i0zFRWRpADimKDXH6zCbPcLfFfGRGRD2ZbbY8LRbY4zknu59xND2i99
44VPL6ma1RIMHGRXxzdHuY07ezgzUttynPqC7vW0SgLGD5YoCSrcn+sXnBibmTEw
HY970zeur3zGTebxwmycMNwj3NJx2eUX/j2fBnqAqlJUQq+4JmJ1tbOuzxBm8Cho
EakL6K7FKNwkVvz6n/1C2mj9hLPHCzMHyruLE0GavqAUzXy5XhbkAQ1C1kYWkCU7
cwn+RIW3M6jxVqUIzOdpGDVL93PVO39Y92lmAMsjxDM8SEICUZrJPgNYqPvidi6F
V0bj8HrLVY0yl7ZD+wnQWBc/5hxD43O6yW5N29JYxjTGHsuocYvIhmQDpcFLkgDj
jRqKgknQuczUtzZ2CLVdp0R8JM3txvdiGaRKBzMTxp1q7Dc+WCl64QNiO+N4DkzF
EWEGtx/7NZzfJQyVigpvpRv0KVvmWmHRrHE7T99fkwYLztLQiov+Jcg9SjN6kgRN
oIa4LbiaDJ5Izo1SW4Vnm5uNVqvdGvI+bvf5iTGRhMUejrBSgWAV3yWeogsed4Gc
Sjt4aFztlVLa1WeZmHHXXkgUpJtfWwCVB/cgnjU+P8st+VW9QIOX+GEpadKI6xqG
1yaHHyQf9cTuuvnTLGHXeCiLi3aexuVxRzi0f4vxbkpCItcp99sgB1Xfg4HpsfWr
/vTlevkt4Bmk59f2Nk4J3nsxcgUj/nufzWyKHCcR5zoWJhui8ILaEh35d+02yJ90
p/TeCvL0rEq67FIjA1FW9usd6z8liYH64lMjan1hZrKOl2sRStgUFXTYpqHcArPI
pwkah6q9Jbo0h+yUvAv/nzLowZPsw6yK5OqqcUILeAF8WNmmgrzOuJAXg3QzwlU5
N0hi2Qm4KWHOFF7QbTNuIS5a7Vju8q0/jumdTjgJLktyHY+Mm+TK4XtVRrvAJOBE
Tdas5B9tJHIoxwCpD8gHIPND1NQNymTvCRMIEctCG1uT+Gwdy2J2+QunO57wstVa
sGO6F88Pu0+NblQOlV7/2J85aC1T5mW66lKPumN2HgCs9FiGxFHO8E5MincvjNeo
qGG1ZuVZrkH4e+oFkxDN0WFqh8bSQsxOhZLsJZojF8aJzaqkubo23fu623DtGTlo
teOj427aGOzguELf6qSuWMDOzqBHK9wjG88reJdxr2FVzvmrwOPO6YNlVvT/qRw1
jV/GhpSvI4hWXxStK4cD3IYraio6kTU8Z6IONXNJnJavr9BWov8B4aVdZMHbLr7g
RN+6ATa7uOSvhxri4sfW1FZAE7a06INk2sZfqWZ12UrY/RXLt2l4/9lgBal0pv1q
zPnopFOmMrbrAxQXZt1crOxGS8SDSWzjf0YALAIRnlnWiyVfOuPoIMoTvB7bOSBT
8+bAkHU2xhzHdvbykKR2Me4u+cEkfxqdajteXn5WluAxxraSimAPiCeLfxdfbtxM
Ljw8VqEgZ1PVB+6yZuK/97L+uBZw0DCqQV1KKku84qFuQ4o1OFhNfjDNm13Ca5aa
JK5TrHKrZbQg1s6Pmu11Pzeg0G4bIab/Y5s6QeLAP6H91/BqFOh4WT97o6d66kR2
yN93DzB1GtqMbgzW8CdP3Cq3zcjaJLjX9/2GIWJfxG8tV4+SXvEnbCYNuD/boJJf
XG+QQHIFNEPUAeHLAY/0Pn3ZvGtE7eYPGXtlzz+wTdY8Mfcxoe2rLkl75XnKCh8b
ufWwOHvDJmTA5WUJ3uTTBo7v3qb/ypIf40j+JzYwRmCpdVy3Abx9OvLtUTWZgrqs
ZxDsPZoZttJ947kwuvCh7DftCvR5FAyIpmVov/bgpb40X26EJZpqf0/qFoQkGwHa
Xef8Ud/zC4qUkgso7VrtKhepxKrX6mOZikWgWFCy+hFyp3Qo4A6+Qe4/HrVbZx3A
muxMTGmJeMV/RidrtL62DTF30A2qIhiFJu5zaT9SQjkDgadUaNIbJ2DLegNUDw6X
FoIhCXMoblcbYBWjju59MnX2wT4FtJPDUMeOSDMTjvdU4c7cuVxmQpAK/3PTeTWc
z+QTnzEqPirHELzl1Uci5igJJCOb0esExUTQSb9pnDUrYBvcdinL/CHuQWV72Fi4
QzX6ReyAVg6yNafdrmN7eF+7C5FYXOC90W/yuJQ8dz3tHQaqUiBgjIA57dHvDyQZ
3PUAvVbykT/04cYClEhhr5xuF9zEa0KtivYeYqTfP70PE1LEcaKMVWx38/shOdKQ
HfVbw5EIFy3Yz2RjZFIOUxM0+CGZNqXo+/OSz4P/mpjbleaFLrhRCit69WQ01fS7
MORTVv6jkNQGAhl1Qn6c+mdLDDy0yLI0AOfcNCnt+NBJZdykfvO3mpwy9k1T8b+1
tYiZWmvudBx3rC3yqL5iDL7I72JZ2pCAg1U/GYaFGr9uV4E9Fdm8h2PJKvnvgK9Q
IhzzNOVFZkiGdME3IVZKSvORZXgPZtB4N5BQkPLwNOkG0+prqbngzWNhIjOmEKSW
1hqk40t7IO10RMSC+JAzXppfck/B0FG93LGl+f7iB5EgkxQxqbB/95itQDDVXJSl
kjYyqfqGzNW2Qr2W6C272RZymHXq/vOflkF1OazZPoSZACxrMN3maZWL8PFG7nGC
aFP0FSo1nGFdVbwtQmVNvmSGkqUrzyoY0U73W7rB05LXloq4KTACBMLgpAyXJlZo
2d2S6QIse1kWLRmtNlQpBMoP+vWe2l0wvqPNjAPQARhqwA+SrtOPNM1xIDwG+omF
yYt0F0RWl+BqoxXwNDARLrsD8tYinEffiokL8DNUECWGbo4PFNf8Mg5F5MTonv4E
uEFS96F1YTxocUB4dbSkB6H/fpJtX3VYP82Hl9aiu2ZrBH9OxrUZDF5+1Mc1aKe3
xKvmdtqjmD/V+xwj6ytSyIgDirUVfjqG90N3zG+RFEIPEFHaHdHBC2KYPaLkINkv
PgF6enDkmQV+NPS+EgaeBn4sORjzR+qr+rNS6MamJttcxqnUdMhxN3ZRYOjEc8ET
QNWrVl4ITZicHuqORMixfr7dMvQetSlANVYe+SLTxuJG0n2W7VPwlGGhYOHXCUWz
0u+Zj7id+XKcVYGosqkOM4NyOrtf0JaTFHSxAGoeItDuwvLkah5qSlXzOCMgvCMi
meggH8Nn/Argoo/DR0qHUmXFfUtxQEnbpidGBcxkPiW0648MCoAeKuqVL2muLvK4
WGUIPXqhO9zLS6R1fpqmw3c7o2qvfvdmlmFuY1A+KF6T+kfeeZMa72x9/KwFvdzI
zvYQOkXfLGZ4eJ/9+oupcne4kqKUYYSg/1xiHwaVVYftlvjrC8b7C9ibjL8PpEwO
OCuDzpd09Mji1QqNP4T+ajbS74uub/jWL0GrRedJ5aGQY2jaOvSPU0Th/ynyHsQQ
cKHg/B8iEIWnCoPi49IN08u7mNGRpV8o5aI8u/T2jZ0HtuTeH/KtpVRKm0KCQhVh
/P6Hjsk3P4yUFLqQY4aaNm5i93toGFOweTD/lZL0gh5p1KLC+AOTgXK/KxjQ5V+p
rq9chFYy73vWQiUuebhlw46+zUl9lew8e72Mf8x1Br1QckAoxCHq4Vprd8pIeNy+
gTgbPJWNr3EOfFGhMxx/ROxBBF72Ri14DXLLxyL10SSOKWAYlEik8UH2/uoCAhAO
rzgRvrpiSFni79dAaNPRZgD9QqSwsSscOqUtMmRfCdw9fH9x6l58eIun5F1SlAqv
Vr3/Abs0COHbb1892IsdT2Nayip3jj9w3glwB29/R1+OwLHO7nIq+CCNGy9Md54N
Ya6n5oaZhX1p+ywCMRmuLkG5Jhk2pdQ3Jh9VvGUset0/QiFpCniHpxBp6saiz2ww
Er0z2u7AmilHJwb7N9d/tVENJrz5lIVhgpqoFH9D+5Dg9rhb21bVH6oNnxVHm+B5
YJywGmWDj5J4gNE3pOP0Qen/JIzsMKaCgU1rUg09WnAbpGRhjma7PeP+8b90nfmc
R12bnqFUaSM1xlPLDM1vlwrPP6iBjplVbYrGKWb0gx0EZavzcd6cEedDz7uSb8tB
jYYWul19KqP9NJxUbKvv3zhPBM3YZaOsQHQw/mohF+TjOlbkGkSHWplqlFroqxGr
fqsKW8sJfK+Rreg327efMYZgxBp5IaPX5Fg2D9jDlMkyz7jfAj+fqRVL+yf3ea/m
RafQnqDsn1YoamRnLkletKvM6F8SHuOLAjIK4rKkzblKhz1HGT30fmObHetlVpi3
/Gtg3/Omg0ys9ovjGdgHOdpUTZSwQt2P6L6uh3o4UT8cWfTZdgzGEzJv/WJi5Y6S
G3pX1sJvirc8IMqpULDnxeXtSnsuRbVVY8EYLOsRbQ+DXI2JAjatd3fNZ4Ql5mb5
DWcM8M5vasc5PGHJTL7JGk9Dfv5Pk99xwg3ttYETwSzKkfa7rP0JoNYqNyxaWQkk
mGrxj9NlF9UTGaK+gbrNKX8lVO8f2qroRhK62H86ilKLJ4kxZSA2o67j1UNadrAn
SelGDqN4y6O1HEex+UdyNpgQSQXULGi+lkndVj5yVWrN6GcluYPXKTgvnRWHXPzg
sr+IyJqojm0Zs6YL9bcfeAnfyDnr2nd1WTbq/GcKeDnhSt8nw6t+oyDVdmTfrUTf
6PjvYN/cv9LDLMxoTN8YH7gEMhRyjnhZD8HNtPtDH8E+ibSnLJ4BiksiOh71MsQm
lXmhcZlVrlHegUI8MX/HCA2ufegtUOuvREk92bhnQmffuJPGxdQkDkpV0aNbo52c
RZW0enqATy6CxD/bg/0LnQXiD/Q0yB6+De2BQU/U6WTPWwTSg0QwTqC/UIxfUlOE
7jObZUghqEG56sjPuohZaOZY1kCFqRoM6Sky4ZT/AE29FpC8kjdJK1Nmxke4PCKS
ULU6QII0m+3gS4diEoexNtZ4B1Pxj0zUfQJevzczEfPW+SmIN79cMQpexTeTlW21
cFb4R5rPXl7A7SFPgQliSZd1Q4pBVfpURacPRQphInkIxUHG9t7oLJTBNJVwk+lI
/UHME77sh1pagAa3he8Ab05Uk6Yx+M+ySGs8CNhqbEUpqCQAFfA5QbsKfCj9A9v+
dGgEGz04LukaSQ3oL/ixzr4JNwTzUdzp250XmBYJ3+0jL6Pi6mi3/pwH/ZvUl9B8
qGmaP0PhxjSZ4cPko7O5RIpLNNpZaRmMjXdE+yz3XBMQlMtFpUw05dreGWelWLth
KPRYUk72MQdnhjSdNCToP5aDTKOtm1G39G15PQFgJS4YH7eFShMpukgRjeVrvpDY
uSCjv9oxMpAhCoTeMBzLvwF3Sc/maUTrU07VKmOun3yJpZ4DA6cp28VDWv6Vqofq
LctNxbgwG6prM8jS31/+RuFdTKsirpB4x5RQ+EQMCVekh54iouwZdTX8UUZKUMwh
6fVSdpHbKnP6aNKUiwxTDdnJ4kKr2dX6eInTQLqBO/vf+bv8nsYp1D4ZnqE76KRF
5woju0Ph3uIHzsWvJLxnIWcWIo2VOqARAn7qBhcaETHUUZh3vItR1wsiSnrCIlce
0HTU4mcg5EesCukn25AJRhzgdtNoM2W3AGlXb8i9FC5hs8Tzraoc+Mh7tnFFGQ70
CmSUMl/7rGMciun8JrDZLq8rJ2WevEEfB8b2Y1sty3p3QIz58kQpn80KIhDdFKYU
pBoaPFPs2NegJhwnAdjGotJrk4Lqd5QUB6IDvhh+J/9YyiBZWQndo0iBl8K8ncYz
VgXEAxgYR2U2iBbh+bF0074uzJQS4QBE5DtCgiedBY6jywPlVQWy695m8fBnPdOg
ZXy8uRwkIemzbcgToun0bb0f9oYyFdO2DkPimUmxF5cxryzEzQ6liqXBo7eQ+GOY
KmFevO+s88PFVcLOOZQ3Z08VhQw1WIL9Hx3gDFidgQzdxbqHMhy9P8yt2WKYJGab
3RoRN2xH70hU1sM+uP7V8XRDf2Q9LvoDbOAq8XSaJFqfotFTeYJ/Yq+Cm3d2WtRD
PkkbASCdZPU41/T5/0aJY93efQ3zHVgMCNnKm2ZOHEz1NI31SY8seYZOk/JTZxcq
kOl7+bh0v+vDZ2DkuRYBGwGR/wRKBfsZs4qDzE1Dg9XRedmkYzFDy7kDyfVutaHl
IIscFOh6cZexMN4QSJaUc2TqtRe7Ulo3uvbAq3yIbOn4WZjy3gyPqzM9IVW1O7nF
zBGNiYc8fM5H2u3IoHNrIulBbYv2hjEmf8GhQ4qIPX2XBV0+SLQE8SeY6TSYc0py
siUCZCPZ7B1xVY7vOVpou58nbIuWEi2EoCdwWgTmkP+f9uERXXCvJam3oRX03N49
Dbd/tdbxG1nARTAj3eOTi09SctUSkbQU3e/fEbXY4gzAPZskS12JvHkw1XqSa/8z
faehoahbrcyZM1jYPjg2LeY77LVRIPFg86E5C18Bk3GXxf9iiZg0OZDxw8X9IgPr
n9oavD398GMkxAcKzmIHpTuoOrceAXHbg24BhBzIDAdsX0jbr23DFVIwfODvr8Pd
lfwY7DzJoxBOhHOnwC+6nq3MPQ1g+Vggud91gCLkFMQBVuvVlVk4yAKMYvXVqZ54
c3SljYNBca5/RnuL5byDiLk/0fmzZaEbJwtAqCaaZH08uz5Xm+5MY5xP8Kqvr5EQ
kzAl01bQw1DS14N3KAlJ/iCpBqjjlvd1Fi8XuaTbaPqD8VL9vAZL+/EargDZNcJQ
qeWIAYpWFdWFRfnLkgSjfl/Eu4k/an3yC2TwthPWZ43MbKdp1jNPsViP0QJ4Y0gu
f43fAZSXMLIjbAOFsCtY45ZbiJAHRt9tWfAWKmbuqn8Jnvn15vfvh5spaQUu1xXY
TjdIwe5B5BFTApkNLw2+FgFvIk74mGpEG+Z5JNQuGyt3tLF1HTPGI/9eH2Vx/vqz
uQCQjtuY4FRODbTpkbL6mjjsfc9Di9aRM4yebLXHGKbN5a9SC+nKftiPICuGyvG+
RUYlmy8Gk52UCeBrsEzb4yN6s2V5OESloe9Ryirj47s3293IAje3iki1lWVzjrbq
c9VJYEzplAoyYyUFe/fJ7pDPFAxKdVhL52AUy9AUvX2uj5x/eQRS3SrO92QYtSlj
SZV8e42ayo2TlgczEssndMpSIICGKRI1sNPzCLMAHSOptoQpOqOtZc9iEa+cAPja
cexKQi2TxuWfeuV91MWX7QN3dBAq3bDwvlGhLvnzXiQPZonFRHy/Lde+FUjlg0Mf
+E5S+mB8Eawy6H2EYZXtYf8dv6mZIHkc1bNREm+sKfWh2cFelUx1IsSoVDWlZylT
24nhckSfDsPBCPf8hGMOciVNxswOaFzo1Hxx/xAzhATOY1Dpebz5cxf3Fq/qnZfH
bcEc0dhSg4i8YFSNpr/NsPYtvAOlPOwe3O6PUVisGM7CR/NO6fDjo6oUpyDxPfXa
6OUe2Av6NhGv29H68KOy0gAh2Yx8pVJO9hxXsQirSqZetdhzkI5v1pHuer0zH8eZ
0VOgh1nJkrSHVb3vTjn1ZffYGQAMSI4WYOa1baKTES5vgGXfJ4ZtphavE1n20GNS
UtftW7ZdxrhqiGbApqQ2dzffWYvJBwPgsCcJ/rDOnWlDdt3AJ2FU7IkfU521gD5s
qb/0LDXaL+ldWHGPIQAOhgpU1PiaKW+4vlymJHV52iA8o5+j/0LCyZGpfOzttuC1
adnx+aiRN7yeMUEd4Gw1s2uNQtcr0ld3XAKXbNmTC3hotq+ePAIfU1s4PFSbZKv1
Q4/U82VHqd616kdT8RducBADYo2ZM6CpF4INv7+g5LRMHCx9JXf1iq8v7zbmjXAI
Thh/2m5sMpESNACNsHQTRA9a3RsHGCs6WkpTWOGCUWZh5GrA/IhwgB60mSaiE0EI
fTlZpqzK90qEUDCYR6txkLI9SUnxSEyJ9FesKCnxJJNtBZHmNgmWU5jb5hgnTpAs
ihiD3cl+/EpO1Da4UliiUV35QkTVCc2sbHTjueiHzQtgQ/8dQfWZIZ3I7eeHsYBu
lUbzPtukE02AlFUPwAnsYlyhgCuDpLUJEfvkL7reanXDjbCq2C+QgCJYWbdjqrLl
J4i4QaECnCNZm6va2S2GfnD0tN9KktEZ9weSmvsHD1FLHFBdKKD+3TfsHA3Xb3e8
NjbhqLA8M5k162VgcXRW0Fz5uNt8Z9QT0sqrymJu7454K+YlAJOT1RVjqUe2uR0S
L78miMSFAeXono6UT7SpZpSnhT2CGuMD8zZykDwtO36V8h/JiEuiurL3BMQwJRRN
Uq8O6GqwfwNwllKxc+nYY8sl30dNDJ6CxwMR9IvjMS9aYvBBetdHA2y1ZVbSiWSr
rG0YszWInLfTlhPEXarvog1tChBSjpuY2mhPVPj217wd0wHoy0R6I/uil/D7ThPl
DRWxEXeOJEOMYqce1xRlVuLIQyU/Am/eSBukXjTxcCkqMaI9Od3LTL+jXE07VQ7m
pMWKo/ebZvM4QMdzGGxkXYgmx0RntyGLtkEcyTX+ppedxwYkz5c1f51arX8G8BfR
JajXhDN3EpuD1fn3914CMcOpIaS07TOqn6v6ulgDt9xHvliqYhLBuNFKEF56+Z5u
l1R+rA4Rl9oZTuT5ppoRpEQ9T2cDED0iD3fEBkTZ2IizuzXrI/Ml9k7UPJ6LtWD2
SdLYJ6y8fGC7/suKPuip+JEPxCcjGZ2FBNrAJjD6Wd6ef+lXPK57rtJBNgqxCrQc
4NTJcFTpKb8I+YMydnMv/yFOGsK3+QI8f7A8whJJtsrIGcGwCSspCCduN5ZQWwxu
DJGry8l3QRebNqimyeoOhHViKhWiVQIoH1mTnLzur5kYOI9uA4HzKyC8Dk1XJ7vy
gpFPIBdCc2Vgk9JpYngGI8Ip5/BFpp/Y2G5vuayKWEsXkKq1xaVZbyOokoxF+Xnz
fBORfwalobvbYFD5rE+iK4sJtm56ioOCmPnxWxv+xhUbMhM9bfh5gI8/DL6n5f0B
kI6HCTdSED9MjlydtdHt9GvJgXe2DOCuGql9mqhvo975nzjrsJ67J/UpC8zf4TRV
oI/6iIHtYf6BMXmkX10yFiOe0Jv6r4deNG0tF4C7TkyePHYNvKGChjc9J1vM4M0Z
qBG3HN2bMcqV40VoIh2m9Cd26QkGVkFXdIJTlZjxcGWGF5BghCu986vDhI3TPADF
VBErXWyM+P/6lfo3q/M4oDVlZdkciUJI97hC1R1tYFEnAUQxLIgNUYVjwwhAbN+e
e2BlSonx/UZNfJObRnBtbL9gBB6MM+hVDQ9YaaKJGPSOm82CCHLffuijW67DVPfk
Qy4M1Hi6bHaHE79HugQ5XrMV6fIBwX6HFnY8l04Y3XRdgsoncH0E3dRZCZ+39Q3n
781ysdWKFRj3I0Cxd2rwSDAN207zHGtwu0zsfESEmiR0x3r8N1xzNccaaxf9MBPk
96VeIdNBpfNK4FpP3JmknPrjadavw27BDET7NHlJbT3+aYKf9f/V0MmiXHFx88gy
rOz6QrJh803MBQrLa0USVJbmxh1744QKRMgrLLzreJzcpd1MWEVnhjjIbtvuD+cI
dH9ywJBo6IooqNugW4XqFVP+SREPkXWeGu8sKwa57+VWh+SDqIZS1HM53/gPoNEu
sacmtVmcJr3vwA9cg7hBGecfugYGJlwSSwl4FKJah6Gwrz6rOtje28w9y1Km+P7u
NJ86+wJFIGFNxaG9PctVhFkqgJT/ldeTR9mne5XfKGH5pFLXXQM/5/EkVj2CKf98
yUs0r61TnksoWNzNJYupNCB35gmbqs0XjHfXjHczldcLWrWsn2P0O/y23tFHJeBF
zCoempDEGq6K4bxY5jYr9Zn+Q20Jy+jwORywDS6u8Ub/fLnFtyv13guMhYXKZM3b
AnGDhc7nLYjot7/6XbsnZ7FeukZiXQmJgaZDuOrfgHGpInqZMFEkPoru/YcI73MB
K7dl5DdIZ+5hcJCAJ3fMl/kHDXf/INLR6RjxyAbZnpWQL2UiC9PtVnJR2k43tATO
BJneJBsyM/3o8t0uyc6o1R7fODysEdXFST+PSLuHbtlN2/Fu/5yYpE7JdYaWzml3
SJ9l+ApziuGis3cL6WEAv3vLdEbUT+1Enkf9Rg1MtaW1UyG/RFYHPS0blnHWzvUW
fC6rDql9zetdvf/i3tAHqeC2gY/8cH0PN+irFHeo+DHgGibBSJCyPOBLQvKwaY+N
W8YZ1tRDmgFYMBbY6uZZulLyn24q8Yor3luWocBaex8p9tNvg9aY+ZjBCIhB1QNN
f5kEz8V2oPA83T157KNn/r8DdgvO4QpHeePIH/+O3K45vX0dZBCw24uoVtEx/b7F
NQwu+l0aktuW6g5zUT3TtaeXs5IE/6rv/BCqkMY3HXHLje/zKsjxjw7WwtO9wO49
23W36U1fo1JyUnPxapiYExqGXRQMd20psnV0/dOddBlZCeKnksb4fneFDJcR+BVe
xqZFgMQIUjsH6qXsc+IE3jmVkV7zZtfREuCTskz1Qy4EfeG4nhZy50jxoL6nWltG
+/Z58yg+NtVjTLZRq+mogBWvHCtbOCPBCRymVAsocZXrXI5UacdS1pMyUhg+08+y
JUEfImjL7JZLohVPwu6WixHdOsS/IqMMOoyGWv5DuI1JQ/Ipy8p2CFX4ugS8uQph
Na6gjVZOgNqGz8WYnL6ccgOMC+p5UxH+JfuEHagQO2p3od79Z1fC7dbe0E4qD1PS
UkqSu5b1HfEqfvMvp3YR0VMSEMRNC+C68X2eTs/IvyqDRI1cSJPrmOJ8bu2oYfmI
c7+HcYzJY+Z+I7pUCJEHaq1GXg2Ja98VbKQCCA+KIV44c6p/nKON2YCmp/qjysuS
3ORs/1Cw2yJE1b6kubE6+GJU07Na3oQJoxuO42m7mc0/vZBSr3qkvA2UueaG0bdK
7IvrwntqsVTRMpSjQBpDERelkFJz6MSi4bgPOokqPHfWZmYFrW1PzjrQZTGA/h73
Y1oAGEQpmif0yxWdtzsppgqM9FghEGSAl6uU0xZnKK3RoQ8VHvGktOMzZID874GB
6zLgBmwF4rD1Rc7LmnnnbSipM+8Psj60Z443yqDzXkrPaDRoxtNbc30QOqFSRe58
0u/C1O78hwVuztCe3RSy9FKENPcc7jhlI9KdEQuMOG9YffsGHoxgjKq7YnHnyk5r
aY3nKdjEUgqHJhJhGhs0KWGB3QbkUj1vGTzBPh++zpe1gkmOxb4U/w1WLsH2NVJz
3qiAVKFE5UHvNksB06WseFmqlpxRzOvWDfgM2UauPRtanbf6XXcrtdp2gRJTuby/
oSzJ3818+gsbxXYqDZMa71s2HbUuQLwV2TXG2Gp5ssWkZtXIfN5YIMuLhKmh/zK4
r2XRd4nIVdsrrOWAllIW4KSH1EsMFXs6QDh63YUXn112izkbGhhfjxLFEo3vaoUX
CnH+huY1YW7/mFxoDPajDc8WC8M+jy82xe26kvR43N9zSmhRlhMwVC0nbjpwBZWY
T1HF/sYiiXvzcEtxSoSnZ0dH4nzKCmNC40c8HCxh8Ip9OVYCebJ3Lo7bw4hbpe9z
qLnaSXk/V0rdEnftB3NVnW6FQ5+rkNoiqJVolJxhxrOfZY8wI1HvaTUzLwV7oyFp
L3PXgZ1FE2m3JigbGVoCEuDjOLJHDMARP0NCZPAl6F4HcgIYcuGh7s8P9RR3A5/K
Med6D+qxFsC1mOhdDxvf/6kHod43AnMLBRh9A2/sW2L/Le5tsDIV5TH987ZANFOQ
hKJ742wsru/vJ7PWDmmocv6YExKQdoHxNXW+Bycj4STlmw8u7bQLhSrAs4hNsnbg
z5n4AlGPy9V+0AB39jewNHh1I8551jD+Y2VJbD/ysnmkvgRb7GWLyi372wNHgoZK
ygb4FM2vmXM6bxHAly/b42SUsaFaCbp2LVv1JHVLLto1VyRgBrbU+AVKBE9/NU1H
LQ+PxHahRpsap1dCxvcnOQ7Ba8anFZIuvHv+pI7I6Q4pFvw6ovHR7yLc50G15SKT
eAcC4Iws6nIYI9qeDj5/lsNTZ7GD8PZhdUaeRVDf2Mm/Hcqe0WursIQznh4zORHX
zLQdUhuAlI/eyuIrVV0hBnnFw1lbNnFaquLKEOZmE5iPax7iZszonigC/66tsh3k
QphpwWB6kVSKNj75zWND4r+TiwECO2a67LAPMRmTfdD9FtgDZt5pJBIIh2w8RjdZ
kxar1OuUlbGNlQiVypJlkatQcC0ze1N8CrOd8+Nqi+IwJULADKsW4FMZ3wUgJgZr
qHh57b2H+daJBgd2NJB1MXng8LUZcxxW7fZeBidzPxSLGrEDP0aAtz63WQOgnlIZ
jmBl47TLYVVOTExCqK1E/DU6XZXECuLevklIcI4fH/14Xd2PNOrsMSymO7k4xgDp
aASuaeK48TvyOzjQnRXyFGqoChGwHLkMZsXAncSjNkWNzxDVZCibyI15b4Hud1e+
xw4LZ+OvhTfUFUbS9uYgZOUaXJPJQV1pmG8BWLoZnapJ9j5Omrkz+bK6qwxKUtM1
m6iPJ30qMCa90SB10N4djGbM1/NUEcugB13rnZFk7xalfftl4DuAr1aB6EUsNgFw
4l+suDKv2cTtXfPnx/zSG7wlMY/u6qWAN3NLnPlSnuj8QFRuXwLcPOLKaAuSpnMB
sCspQ1w4jpxEkgRi3V/SOTaP/O3rVwXue6BI7a7tikuSLbxjSFaJiVdUrSYQcAJB
OrXIpzpM4wb4Y0cJjKqzmx6aagOxoyFdpboAe7rsYJno0CBg1MH/rXrBQtaTvVFM
9UJOG0nKf+81Yh4GUBK0vAHnX3nDtmE0zk8tEzHGL2HV5HvA88QEv37sy61VI/rh
RnMf/f6rAw2Kjmirzm1jOZZvP9kaCOxovOz8gYf3fUPsOwLDaJMRWJrWCz/3emDq
LO4GAdcPPqUkupzPSnvi/KHeNGa7RFbixmLnQ9O+2zI1R8Jes5HKTADIvJMtKEzm
tF3JHt+38iAksjbZHTu3QtT9KQsVumbTAthQy9dXK5nDHx46kIp+uKNSvmPjeCgP
0Mm515zuhIJ+alFVXUT4+um9qdTrpz3yH4Bvq/oHnFtyMnlREEYDfCKYxL41HSsz
eLJHNPisS32sZcicZJ9215y/MDJUGIBpcir/+HnRbvK9ta9Q2D+AM4qx6dj1ojyp
qgnJXj3Go7b8nNG0azu/+c6YUI2ai54oG6n/dgQd/j25YySuW5KQ0hSF+6579x4n
NrZf2nO8FOC4yhOCS0v3MSo7V/29D8Ff4Ck7Y8xe8KettcBVjgI2nxDwvlFTJmQz
EUjmmdjmGHGMswVOJBHcG4sWuqL8jd4nRf5+t5dsDGJB9yqDiNyUjiNu0lk/1YKw
hxm8+amLQxmvrkhf5BROlsn95KQORZTi9d/a4b4iSyydEh8NiEPQo4+1ygcrlHXC
/MQ6HRfhRrns60rhsLB04Pd/TJd2ISmjr0xPYxjkuP3QdS/KEgj74mH9eBU3UAm0
hBQcHINJ59sQbqvkrUD/ziQ0aqtCN5WVLX/sWG0OtrYmR04bZDtxXb2lPwLbEczp
P0pRXzTlCb4SQhQJqYUXZ8EVMCUO3aY8dx2sWODwJTKFcixhMbZBo6FlvBqaPoOK
CCcl4QTz8p3AVPyPnn7i7n/VMA05JmQM38fE9wnXVwlj5UsmWtsfOatBJZU/h0m0
QvndITPAzjSICtuVsKy6Sq5O+MvuJh1npNE7ow0EPRovbmBe0D6GT12QLEhe6m7A
iwjFBUoIXXLV8V4v648YAMltt7gVU6mpU+hL66B2Y1oPo0VzccbxD9Jm6ZTvha8G
rbZULnB0u67GjkgyFQdTaF3M5IhLUZl4VyyndVQ2vdpqZPxzNbEYTvFtnkfdt/3x
01AuRUmZGxAY+fkeicMBf+5BEA/yY+BUtETBXZZOAoVj5tsleFX9zEeFvf+pP2+e
WAZ3i08AqVbc9vtK/aoHV0cHMKwEw5tlgN96kGcKhLyM19gnLOyGdgLxK7dkzTBr
3t+qX/ndPrEZLp6qEdjI8sT/0hjEBlM1CnvlWSkP9mjTzITrXViy76FISY0+aNex
I3YNAq/tH5V29Te3vDe6JhWv0KhYZusXrqGVu/kNcGAtpbYL+aHK5Vg3kCAg7w+i
m9m1Ag6B8AMaL1hYdzqWwA5ffo2/Lq/Ov/BxJj1ihCI9i7iFp6YOXwZPaTk2AoOO
sa9XnqI/Q6CdnRxFgUrMuDy41xBlO6JF5pAWWsvF3vn3xygrlhs9tgBnINKyu3DB
VD34S6NjnJF9z3u7o1dYdb1L0+uREUw1kpKdtF6WucBanKNhnnrSWIZgady/yoXu
L5ZY6Vrh333/6XENWzY8yBe/YiNeD00TsqD9o402l3dq6hNMj3IzVm7P/mTPxF5O
nVUjZ8aJsbSPE7pMa9R5BR7D4idCxIcUt15ktulMKq1/4zpYOqtPborpVbaHHsAJ
sqeqVUEXN0HHg+qAtvDomLg7LoT2zq1tegeZp0ERpeLzX4JIrORQCh5cShguLHrx
8oPNgFUXCZU1K43e7P+DYPSBmUwkLClNAJC+TM5O4IcRQWuhFJrWWg8X7+BYzsBr
ZJtBi9h0Qsf0zUAY1KzQmC0CNbTOZk0TQZ1IMwhsbIIUBd0Shz8B4EmLL55BbyPf
BEj1VfKLohgh7AF2UYX7u8QJrFjx8L8i3e/NpMx+hV/x27WTDWyW0fJVH+JE6LW6
nctOlAYxWQaP0geK7N8wqyNZgYHvsxVQJ0HRhOM9kPFFmLQb6otQLaxDECRDWgA0
5x5THbnZbxuWnAvqXo5z9jN5vDiH/6GS0kOhyDZ1D7M4y14F/eUBZjA6vstMrZAL
1BLKngyQxjaZJXOOV5EzOnEjPJDKlbk+RPFaT9oe2LgU6iBPJsI8A2lyPb61djRr
Vqtnlcf3WpfQ0BStVWR8s6sYZhpudBD/2n14oRL4yQ+fDBoy2G6sKjv7VzeeIWqW
Cr/IXJHP8faSB0hgYRscVkQVBYjPIjooADt1uCnpsWj3dvXGELd4hObTDgj6BDPk
9A6rT6unM37xcD1duhPGz0fZPWoZJR8COwQ8NnIUF1a4TwN1e9GeaS757N+tkrn+
hHo+MHR2oIZo6GEQDhntBdyemGydW45+qaQP1+esMMOZ4b9fVjgqqpEdynLdfLWT
RiSOj5jLzZg/WZmocH2QK+A42WTsOEWm/CcE2LWG8V16CVeELUURRe45v2tje643
JDzHAMMlPTvub6MeYekN59HBci6U2cTPUUUGGsJupJq25+iS6KysYNTq9C5rHKfA
IuP2wpuvb0jECfD/amDVxEu1a5AFAzkDRW3rMO6BTNv40PiXoVcGQ9b5Bpe4Xjaz
TxFyXDO2sEfk4SCn3QLVxLJ6gd+Kqoyt0FTdnms4RI32X1/Xud7QgSXvvQrCrHEz
f0/uvUdL8FCooU7cQkt1s94SQBpEGcrrDJk1iiH9SHWuKGUaM9sq0i4IieEsSDkT
B9yrJ672RlwjCjSO6EhfXq8ueY2fa06kYmulylvovuxcXxiIGHUs7nlPvv9nzxyn
g/lLwDw4zy7/WGbwR/Uy2UEdcQQUGr2Vlftq1MLiMQ3AxiQJAf6/2v7bK/gVipK+
WJRCzAMJMp16qajy065bbIwaICmCEb8MknXJ8CvgzgVbxtFbkEo8NBZeABsfdhix
giz8vR+aRfHlC9j5KxqD0tfiQRL0/8HzF8XsxB7h9erzPC42g83bQ39L4LhXxq9J
jIE9I9GHGDktIQix80gpB1aehoOOvdvh03MZxcuq4Th7ElbpNtOh40cPqz04/yse
ktqDuyOSCbPMfzxXM5PG23D26cFMEy+4AghuCSZVV0r03KmOqufroyISeRn9aISH
2EyEM8oYJF1+TCDCCCeLHltjBO47i61BpDf2NUrH8IbQ+kabhKOoRZ+AGWNl35Mv
C0HuT6Q4KIrT4coXrgjjY18gdFrfdCZM1+dmF80vU2Bygt1GRsHpBLDFfnzwslZa
rb9uz15tdfMst/PbJZfpt/H266HQNUz5J9JOrI36TTDJ/pON2cmapT4ixBQo2aAx
fNMeBLlQZV5TYuRNEkDlvBSrC9wuLqM0qxp6Qy8jKvSKIlZsqEVk+yL2oMlTS37m
MGMOlyNE7aUZm3NXRMNxEpTaOj1JtVl3bCTg1irN/iY9qaIoivLBQAGKc7C1xGLY
m1Mh1xgFzXEr/NGXwMoXodbw4iug4SwKrQfCBB1tOC9IQMudMaW4MO1P0DcMtDA8
AGyDOdkS0nOq+5L2LP1x3DT9T36xa8VNphxJUPoCw4NbC0r10IRTDs4hqjzArYRY
ElMmJ5SMjtUeub2Liyps5iIhZQURdYyJf+p2EQdpBDcD7J0dCMwMrQADTGVeGY6A
jxqksFEQdr/85trqSCZtvH+KUN7O4H0zr+8oAYCkJoe0EpGeu4ioBNvxs1CyMVpz
eAtrPRDcAa585q4KxYugZhFaZ6z0fnlHaqS1EOHvbNmZaNSX9ywFQRG7QYSRjV4r
FNSl6OVorR9Hiplb0FTd5PXYO4YKAHNpf6PMnWvDhniuWlugFcHnmDRTmWHlohPN
MJxE9wMv9h19+Uq0MVcgNp/1zRbnbnE8DHV0BqryXn9khCmSk+Em6gdqP+X5/hhK
Isn3fLzplQABWJ0UrxrQEnLHNP5ogp2yMKkisXU5nnIv/8MyiMywS9x4FJ/FJ5pP
o5UZY/N+uApz1ihv1kqoeMYvE1HhQUQstN6R+eN7wH+/oAFxZYyfjLVKdy4PZGjA
XXAA5fqMZRfyCw1iJI2gvLmYB5nRh4iBbIPimDLcjhxMgMGTcne+Pgg6c/KZJh8H
YxsapTCg2CF6era7SQhBCpDepyDP6VzqIsqxnz3M9U3CA+9sR8abvH+aInQH1pK8
E8CB3/Y3IolD6h2P3siGBt9wi3L0LTPneOrw4utMAoTEx2+8yO8V+OsDT4/wttWQ
yanbBDBM8MPSkeubQzp1oorE1tkIBkx9RyZYD+egjuurpgehe2k9P9XqXa01toyL
eVQuYZC6wW/ZNLbAA/wwsCpVZYKDclZIA8LXxeSiOdeEKsyaMPdpRfKjMsJ3hnZf
O2sOPtLAe7kzOnoDspeIRY1YojWS3nFaOz6pT1jj+eRDfAzqywQxq1XkbivaW4FB
ooMn20VL5wcGtbwHyFaEiH+40LGpUkJBtN9+jglqO2FAvFmNt+cN8a/u6mpyt6uK
Pn7/ajSi/z5334UtGS1dR5/oC5+jgca6No0+2PnRIse90HGmicIq3Daz9KaDGElR
i+liXVbwaiJu1M+1TWQSZcOTLp46ndF0mZ95WQc4c8V/3jDa11SwYFXzLn18Ceku
yPZgMUFu9nlS5nncrl4O+Np5tsVUabJMOn7GNnGKW+DQLu8LoRRPh53N7buSCVtn
3pTMN9/x3Y35Y/6DeSH2miGOgEkYvDGZjCeQno2kAMdiYorEOlBw5Tcp2He1jCBs
g2gmQnyqBg9X4lNl0khZLhZufp9jc0K8iq/2Np1ngSZjDfkz3RtlrwjWbzQLXasZ
0+nUuNAdfJiHs/dG1NTNE2NCB4kq4FDEWJEbhjuA+x39P2UM69MxBCpmcMIdYT3i
x8st+ufzPacRhqmGPfZHvzIiHsdel2W1KOb3kU2GW+5I6ytYQCOsN7KsqRLtKr1T
DfakmzH2XQYb5BVmvCLBbbIFHVbcjTP2Ue/yzPL0GoJMxY6C44ZQODGd3cNU0mT0
PeLAPGhIO+5M3XaQbaoBpAVQNe0MtjDtdMcovWTQQ8T4BvEcMtd4KtfbuqSoH/Rf
ihyLhwT+1x58sKvSrFkOBNRqDfZNFjBrujEYyzoj6AuQqEXBuI3nN4tKgkz1PK+c
IrRmYVuyJa1Nlkx2tXDdwDLdSIMzeSWvLs8lRkanhbxISVnfYOoejUhAD820PAa5
53j8NQYrYKe3tnC81rEB4siEz3yFH1azn85kXqqHWuDV92mEi5mUsW+NdIG3w/zI
RVKcSxyCjCarD2MYStZ1XImNOe4UaZ0MXmRNtL10J8LrxjqEgDmLRvpjmtvr86I3
yLvExxtv3+ZJcjLtumwMsjBRb1GAF3Wrln3cDgm+qj91JPb4BWKDKi579uZnWzK0
SOlGs256J8kal/F5OM4ZNu/ZozwVQFWDtkoo+V2v2G69HVNg1NkAsa0qw6j9gLN5
PTknUoju1Pe+VjAH+DhKt3Iy+xpTQ2z/sycg9fwLOQuWwE/zHvMJtprQ83vLO6Ej
FcyoMO9AqHGhWezARrExlwWTr2kLLffUsmPSzkRl8snJlJL82UhB72rnQS7xRYlz
Ym31n95bnQDwwQuy3dQ1koQpocXXYzps5q+bM8eLIcA1NI6c1m02cbAEU3tbsylQ
Tqnqtefw/XsY+3VEKdfRDejTdqzFt142fDYy6Zul1PgLu2kysBffeTI1wkD25iEG
PskIFQkeiBca5uXDtbIMTGLb98QSiiYPnef1xANVqtjOJvc9BaNnSE3t3tTv+rq1
9tFHrFEf6yVcCgIDt4wPbrulBqfyMDn7zuWH6TgzrTsGKbB35OOuxeZ5UCZkWHHf
GEhjRCG/ExIbJiCgO9t1FxM/YFJiXKNpVgaYQqa8HYzfj9LPJi8JYcV1e983evPo
fnbJKwdiZvETwUbSyNrnPQYEu9nKzm6fsnhyrJiQEcQutC5oFt4HiD1uwc15KVnL
SKXIO1je9S3EhY+6qufqBJc5WOJ9fUzo1jWPjw19mlmL0t8tYBQWKfyS8vTME85f
EeOf06OoTlCcceQkH4P6IFtNfYGbWm27//h/CyOape0YrV7ZV1EEHdq0PQ3wTRZE
iLl5jGGeOEeh5HFdfuR3qqsxYtgEtXAzeIlEypIAuYvCpIVh5i27320x11wWG62K
HxbVb+OrcFouWPsi86TmSC9xR4wX75EhgwuFkSmbsvpL/ntgPKIJF4zg1c1Ug2Ix
yrQKE3GqzNG6axNKYYzCHqns4VAnuKunus6RAqpD2eMBvw8btpUXlWtOAP8qLuzy
UXwSNpY8J13FAw5cKe73zbZWXuk1nVKQIMX6LZm9ZfYQDKTtjaCJVY8Prmb8S7Gw
pmXxpl4XeQIG1rJaWQV3iPwrlJW72DrGr7pojTtvfZADgFK+hVsAC2zhXQt2nCxa
u3iDuLt2LMr8DuKGREbXAFyj35T8mVE8Xv8Vn4TmWL/b4wFwnLmEJf6VTgnBi+Dz
TeYYRzFLfkdp3vqNJUsmCVNd5HtrXK75djeTirQKNxQlBB804zlsoWJ5QDNyTmKQ
yBpQmEus27cXeKPv1UJDguMDoIJ81chkWSUNBEOL4kjJl+uPr9zMvliUBX4wN2Mx
J/9sLQ5jr3GgDULZadBEczyDus8P5/p4QLL3ocDV1lXrx6BblqPcXUck7rm0Vr+V
Y+5kbmsi7jgEOIJRs0N7jKNz8DAv0vUXihm3qbPf6imv5CZpiCRRINItjeAj+rTT
IYWgobITb2QxJ3w1UIrZlOH760iBJvx7LoH6WzvGn8z06C25XENBndF2Nz12iUX3
V1uuxBm5q2CJEeuqdWgS29SZr1wuVUqFSmw3IN4aj9n3ZuGgib/oloDk8POqqjVH
GzOtBoVYDOC46Z/ZhON2SZAlLdDNq7EysSjvFg8pgSj9cY5SAnCbaphBW9C9+Ihl
vNA8YZmcLV8oqHAszcNxtlfJvpHDYN83KQIGF0kV1Qls7xHcFIrcDe7qRc7icYgv
ZqB0xrd1vHe3p5S6eFbHc8HUAq7sx+Ouwuu2IK36zZXSTkmrwvT2ZN1jLhQUoc8b
XrhNMI28MGO33LKaxlbwmJhc2Rfk3x74vh7sGSBJH7UpgAWSP85r8+xx/QBnCpZb
DKF5sLZQIMnjwpzMX7XzsjA/ZhZsQHbkPbAg3RLal4aKKDckb5K4oDxq29q/hTqb
6CGgxhxfiivN0esaMwQsUW9tDUI/4P2HGq70R0txHuUAQ52rBPHbA3+o39jxGkky
5wOBcAckDottYY6ynYPQVXm9IdSoK8juCOEM/YHDOZe03qTLhSiXXbHnTnh1wkf1
1Aym/y4LC3EYAl8ob6hgo5OtdzeDUXEHh4eOHj5TInY7ssENhoNLIu8p9xQALMSi
kBZe0K1r+PHxUCOzgWcXZdilEinUFPwSHD5MGKXX5VnYpH7lr7eWkhCHuqUK7dn1
vMBkQsU2857FOhC+ObzBRRGl0OPWRR+T/9Q9fy6A87ltnqNd5apV+vT0lPyuhE6I
sxKGQErfrxzveD49+4R1JuYozPjs9Q+TipRxV1jXBvKjAcQKIvMknAJwsuDfbajw
DR56WOY4DeeGrqWymxMiqfvThqahLnEWMUC49J1mHXf9pmQMHYhuUXv7EnxCQxAA
eedN0RLfFt8+frVovbD2GII2ay/gl1esglWwZaMrVwqQNR5R85Ze2wZKKfs1IwI/
4/gV5ieDt8wbsiKvEqUKtaujgZPWJmc+CoEgNotP40nuZC9YEYoHKZT6smtaPENg
tYYIYzvg+XSaAWMGlXWQs/G2rtpPeuSE9a7uujaHwaYwx2H3zjix81mOpSUP+RM0
FVwWEmSvNtnizxtWPRom+MNUhx1l40qZoSD+ZSUBjTHee0CeO37o15kQoPZpUp7P
JqfVj0osViAAYA3PFk5XnPaJSKzGi5lLEM1hQsX/qqyvoS1/Na8DPn3C+odjFQtg
imBhnuyDwxsuYJxIyEdIBjkLfEhoVme9qiNCikuwa8dc/9RorNQRXWy8AZCSqVm4
5PEziLrHewCutPqD6aWHk7nAVD3II+DnoPnnzQdqTI21nuqrnFStt3fF9saulL3G
J2LzVxli+CRfci4zyMmtYxrZ5SNafY7xYp0oEU9zfF8QtMAW+l0klh/6nLhG1T6K
PfbkKAGQyomy+RUXcEiyca7mBcAW0OsNj7Qxer8pNGkPrjGs3leDoX79pnYXsEn/
cKA7cDo0j/7ardrzmuQo7DBD1SBhbSU4peFwo/2am9prkUcWC6dgCoaJcF67FU0+
o7FoXTtDLfrirb4CgtdazH0Z7QGT1NzfmLMviZIKrN/aXUb+WseHvQc0dM6PbEPS
h6X1AgdyfP6vtVJTDh/C67NfilnjTuKnaBjeCwx96CHZAsXEfrFErBUYEWpRmx6R
Fd9bcEPA9S0hecQp5VbUv/NH9sTsCTPPwecqTFi/rTaN2JvLv+SGPfouLNEFb0fr
MVuRfII9MXXASfibMR7PpXL3xIlGmi634641gp/0JjPrrM90X9GrRdqxDc2MZHHJ
W+h10LKk6aruvm6VJ872bir+0bw1bE+SY28XQDDcqcqN2VEpAtx2W47FmA2T37cU
Jkoh0+GBk75ZpFDQ1Y+zDpDgGmhdyfMWofpFscFWO03n7MIor0DmEdN/dqbfcTH3
xVXcfm7cmEm5GOIz3/UP0RlwTffE1RN5u6BY5o2Qqs1m2MI/63mGuPqbdC3V2tTQ
6UyJonSXZtRt9bk2zs2jZ7OD1G2eDfsmEpy6fpn5VD7O1Xp87hoRWJztC80sBJnt
t0qg98bXspCHxNGziewZV7NX8dPLVJomRgyAvmU5PGX6ybwbrN8x+TrYvM3K05h2
rg3qW18uY083fCzR8tQO99X5SQQTzvBpLPqF2Hv5vjzo49tLmxT1f9ViR2QqyEVL
sAqdVsUkcZ7CDPt8A6ioMCwlHKao2Fes9hrlRY9YMgkyfab1WPnWDriI4ar1ppGW
BZYlvCOZZtVz2L4rJF0+tTnq/ovRVrGwmiM+gy5rVXalhmgPvSYZaXqw4VQIVvsF
LR33fjBFrHugoHY20yo/2FJNdmUcfiYKAHLeSBbfEIngepr+YFUvA2tIHmIK8eYW
xfKdRL3Kihxp/ed81H91frEvwggtaCOSzekYNucRnchul4VSvbCIMfISoQp4W9oo
HweUxxywAh/B2FMQwBhMVBnkrxU6rbGhOmXaROlfWqUll1tXx6DtfKqyUaaEKJoy
1M01dbORGJrW/noxraVpDEK8N2KTfvdpv4wi5N4rUEZq5l/dl6NwFNUavlugSyN5
eiFlWO2sMxc9kTD2P0ghTdIqbqFMPbZgWc2qWEIpNKyqB8okJiWPo1zCcew/H+Y9
WCB742b7ZFmKNRajcvdJZjCgpP4Sd/HhNluxYBBDCQ0DnD4K5ePpGh4Z1t5Lsb5O
fSvfrc8t1/VUMfDenxLqvjjMN4dKP7BHP2vC+OzhmF8FlKN8rZuxuJKxgdO3xfbY
2AQeqGBX1ap3hxsmBs9h0+LKcVIrk7FIB6mIRTvRPVzf3zbzmjnZJ+AXdg2rueg9
y3WoqLUdSzUxOm8N+bYZfnW3fwMUevqbVA1q/erFkg6LL1A9puJIjWdxKqFwgpZl
mxdSR+NtnY6oo4zLmzpzkPXWM0FBnoBC759+UUlDwGTfWpERZcx5VqS8xfQM+H15
Kc/7zY33gMc1JOs44eVo4y96q5aWfK3+LnEPVJtJZ9NBU2YDxYLyGvlKiNE/1oXR
YDIT7O4+nGCr5uvBUG2p1pyR//+ToyNWfQbxhpo+POjgCEO0pwuGXrcjDbiFm4BI
bHsJAzabT9SrjiPqX6GLDVgq/PoxMY5VdAdc6lihLPPHKw+H6D4w0O6QkWhOKay+
rXNocQz+/QntsbIQaNJKhQMTrqWWXVigYLn3gAOwT0feMs6qntimB0xtloCp7eUR
RM5xWOX/oK9kkkwIFYT7QZkOjJrSUBihsk0amFmdCp647U49LHVE/89IBpydsblM
Z+0dtdP+X4bE/eK1Lv+B1WcOh5KF5mypPBv9lfC/C7Rg0ev+PUrZF8szHPCozveK
h684uIMHcO4kXKk8G/cPtUDQkDHHYuYpBoU9Eh0kXftEZkegoWLQSP6vtRZrtGKq
7QquhSvrnilpgcU+vNR8NMkvococnxc16hdPH7HPuLOJjdgaozquA1ygekHJFeFm
Kz7HXtH5hXjEjnP0NK/KgQg8ZXjaG+HXJxWKxhJ3xh8UCIAORO8yenGVjm77USt5
8tFAN2zXMtkozEDLuK4/N/UJjkEvxF7YATK4AKkys5P+sfYTfKaMag5/M5oUa8Ww
J5/+MJcEVoNQ+Zt/p/1GTwE2J5Y2ZGYvmaOTx+/nDtAuyITfCnRUtx3Zv8BzypyI
Y+3b6GfBf6ShG8vihN1sYPrPugcGqJ9Qq9sRgialYUNeINauPvHQuwHrNhUZkdwk
`pragma protect end_protected
