// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:55 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gZ7NeEuXjM4/gncUW/+ZgDdL/B6073fz49ZBHyKOc9Uf7LmdBYE7KiSw7HINBmVT
e1OMsvLsCdLex2fO3P6QomNSgSl7+rUGSFy4PjjmBkRp41HkiDLMr3b3vjgaHtG/
ChaU0K/GUnhmFDdGZoCxtc+hbMcut+Uvs+RD+1RD9gE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7296)
1uALYQnH9uW8xmjTW0wo/ANzJ0kBaOa9m4rU1LeS3A7MHVRVPMkutDoqXRMNOt0o
Cnj0HcM+GPoNijRUTPfiLKkF+O8N9GMa+edOo7mvU2OvSUQW1iz5Q+LwOXsI9z+W
p0whYWMrN4kAeZbfUhmiw8gUEiVheR/JeYmPM3QmN0f2QeaQ49pSY9yj3Rvgg6Kc
A5y/2CBSIqIxceY2WXhGEcn2JAEc4uS5J/q05LcNxZAIe6NP6+q2GQ+1qVlYt24k
MBGF080ek7hyxILuZKs6ppOs/X2MqEM0225X1nYtbXhzOmMG4sGbYWlqcKEe5cMu
N/KC0ufkdmuSsAE8x8EhRy0UJymni1Xe9daW9Ft/YEyQtmy1UbqdXQjwaJkBJ7aJ
580/giiTV3iraPun8FASDyrTcRCXn+gWCY692aii/4t/qQVPKnXcW6HQOU+4iM7w
Bg/EuG4BtaXFt+Wx7iHiPW6JDla3ZJAjOdC0ZvDyarm245Org5jvIcexB7zTXZ5M
HkQw6Vb1M6TzHKBrVI2KOGNgPdkAaCB5yv+zV6Hwzcftfb0AoyeMPqblOqoFIosu
boqDzfiN46gJkeI0E/1TojRgKz620VThBLMXgc3wDdSKl5ZaBoUU/bJ40un6Soq8
2iflBawJ8cdDdrcrljhe2NC6U7c4KlQo044cJc5chbjoH1n70CLGkVfbmcGOGjgY
j889q2DcHGjQhKaVsj7FRv9tusxOnt7nPEs64+EJ9znx46NIDSwWP0R7KY+SwZg8
tagfCW/UbSA+9GhYuHfficNCSBiiw/DSctxQ1KkA3akfRUSiJkwjovvDb2/uqLSD
8fnC0UWQTtF/i3dliFDmXY0NIdBjTdHismFMOAtk7CHcBgGVsLWNW4pA0zzT7N/I
NxSf3IctfUbgA0lKz45rPsXx67dot+rUp3Znt1+FEWAVU/gRPk+JdhuOoPLgVylQ
fZyMkn0H+mxzgHQXA633WYujUGe2jD0hpceHbKdRKtvp+D0Ymvuf8+d0EThyUCiN
/Og9W3waUiauChtO2qxkz0uhbdGHRYorDqEX1Ky+r284HJttujGNLARJCaN3gbHb
KAO4Vj9gK9PVxfeFb5j++VjU0LTEfIhQ0Yy+iCneBhXM6LNSiQz8L1UfxB1WyS+l
OoKfnP6qVWAKuN8aAv0ODCI3BQtIFqB9Fo/5BwcY699FCefdFdpe8EeCrEBO5nn1
uUBPBKOnjGdiiZ6MGT0uyPnclC2RIi4uxw4Z/Lmr3tZhHi4967pOvshNIZZ1AuO/
O7EF2NYj0ZN+IZwhqyHY4aHx/srTlznZNbjNDW78Q/cIoT/ktuWTTHjFFIcue2DA
XfVoIUS8S76n9D1/qPijar6AkXeuYGG6UpdUG+BQJQn5QW8y7vIe3rkMpUZ9o7RC
DKTOIC+WrL3p6zfGML7mRHTfTXeCvccefoaVFZA0pWEmeS6oDhVfKyzsYZ2U2Y3l
zF3KIDPl+z6n+ykmmlDBZt7FmyXlDvV+zkBONs9YSlX1UXc6ACWSS5FfLzEMYWSZ
/AB/PEk16Xv5wuFWzHqc78V0njITHurht3F9SI6MXgPddM4oaVFSsd207PzUbV4L
+WluxZXbTkptTYSMfymudPjTfMqYyK1Xev5ROduIXSE70uNmAZC4HXJ3v27yAmWm
izhkIfDzvpMf/lWi84KKH12uR8bmBcUxvF9c790DHOc9R9MaPrGKlx0nbLm4sMCj
PsfN/rE8zK5SK1YQUGWaJfm9loQgXj7nMQiC5i8DUXrc2ThLQpNY2qNoZVgqT24h
AiW6KMV454jreY1SB96Q3P2K7/vwB5nhEja52nzwodx04s1JerORkiIpxoDRxcKI
fF//RyKUDOWRmWKWpzxvnbD2ruKDNgP65rCxy0dGwjh0H+ZvoxG1oW8RM00K8vrA
YgukgQvamvpDjmeiz8n/L8oFRS59+aSh1BgTLfkuyaZ8OjksKyLL+HFKqXmq/nW1
YNeuDCdaan+T1br0xO0JZG3WZaDND33n+V8peCIu1ignTkFuTNf8mnnAn+7BZHQG
OB0+jAp+vUImmCzNynpSbp/lEFK5vyxKS/15ZXAxgMYHqN6oMYSjZcvoJBgyzdYa
LRWoSFObRwDGC+XMwqf2g+hoJog0BXUoYxl8GKYmIcyLIRBe3KVz+u8NYMB4pM9h
abCgT2pxwoCSjjaTdluo08GV2/4H1z0+hJjDvqlNeHrufDPTy6UN590dGutz9WVO
bnYROsX1XPNrJGniV/HTQV4O7QknskII3Iu4kVUZofwGyxztsjODVc2aUhmh48jJ
xtKfCDN3LCjUrHiof2JDPwP627+a8MlykSMuc56FyljZkdkSc1YRvautEfGUpZ39
Yox53CYcAFgiwFnsQNVE5NU85bYeHibekGQ7Qo5Un1gMcUbq8wHL/ZBGdB1k70Id
6gBxOPX0jiJUe6JCBFMQabTkQ87S4Ca8sv/C6gFUqWCqnBTlRyNFHU4bT4fI3v6E
KbV743kwslt04CvaOiw+yomIBLxK0W0AK1rwKPFdwyUk0Q7ejGCkHNte4pkRhNl1
G3qVvpFxDS0/kcOYEGMHIvUUgDM4ECOvn+6xTERZqFCx7ZmvJL1wCNyXUW71T6Ve
ztN+h/s3WBHeP4Ajd3KYtxq9fRYc6ArJCMXNX9YWpzvfcjDlZ2eGbNtFmBLmX64j
6SZqWU97RduF09I7gzuaM1U0iA5z2AtaHFHODbUPJpaocZu+pykZfrf8NOwKSGrT
dtKXrLgk6UJ4I50sFc9Ud0uQb8dh6kWurxAhfDheAUOVX9bqevWIxvjUQ9F6rdAA
ud42fa5LzDNrRt2kmZZU5xeYwDEqpqnjrxg7EeOdt6C9Dy51fEUFGjw1y+aK1wrK
GxbMNgoDCznGTnl4XWj9Oa+PaylhYBDt7u3mZVpXqesLq/C6MQAJW7dSSdfafiCz
e9JoD9L5oD53W9Rd8GD2Z0visKvbzpPPjtasCb9SSQwdJ/dyltU2Hb2Mg3Qx9PuX
WgSXBLOcsMTTPkuepqxWvoZr+vRKybduU21ctNEaAEVIeSXJ87rtzZlN6mjAE3Rz
YmZ8EZdqQxL+h2NYVjgk61VruVGTj1n+fIAiyicJqzpNGp4+r+k4Ft1G2hnebs2n
8fpzPByQAFhf3UHfrPrCUxq+ypnVXhLCGs/iLnNfBSUuW79EyvBi62aTWGqPyCfr
M+1m0N0qPO2ZQlbqUStxqHHWZC+N4pV5+rQEKz3G9SmunAcPGtd8r9FoWHbPdJCp
twkHSpkJaFqkKzYX5nXDX2lPly4tEJjl2zj9kjOLAFmTjnHeQVLrjjGlpIz+OOZi
uiHYbO/uKA813WxJ7W7GSnbocsbQMgjIHzAyjNdn1F0f0uZPvMs115Ynb/PryUc+
lkvGQBnkiuVaVE9P5TsDoZhUcGaPo6viQlUOLExf0FsTQq1SwG8qTFqkVKq0d3nv
Klnitb9/y2cV1QCo8vMUNQGXhu1v9hDZjXKtqqsJs/A6btOY3DXSa6VJoYE+CpwC
d0bXXKcoGQvP1KeI9Nhv9v3HavTNrN5XKn69rdrqQrM8WnQZNruH0YiId4GXLNba
S33qWDHIoiXANHelUNhUfxyejQaWLceRxPNL7NiPC02JAeLFz57y/F8XiT5EOIaS
3kXb445/603RTZn+7W8OIVmhkpwCjaO6qeA4nZCrvwgEs/38DdtLpG5KGwdCVDAO
evmig5Rdhjv4FYSe4hQiEaD97QGIdHaJWGxKgTeCM0l53xhV/43yI9s1Stx4gVt4
4dtucPpylgj6g9Hp4hftUxiRf7IRyo9IOLUj6+rUGPUehCtTWLCF/AKQIZV6dfV2
bq7v7r6obvULT3B2fz3Z2JApiuFuy0onBAW2XKyQkHqqaDaysZAMVvCcwiWPlAfP
ACyGClv57t+nq/R8Wu+VBYbNt8gbLMHPq0ptqXw1nHiP9uAmWmXIPunyVat/iSsA
lzLEOY2/Ur6SKqN2exMofd6ghw6QShiNCR+nDYjziaFWsHEDbX+ZJC9Kmh0iWR8s
xwuJ5Uiy7AaipO6VypHJ7U0BEuMm54mDhV8AYDZ5JqidjCaxThtMHCA86DMwu0i0
/A22JJrcaEpplUbNmXSG27nRckDQNknK2GTgfcbyrP+jBqZ2nBug/sG2jrOp2zZh
66umNpht8Bk4+NBCNzKFkXz5UPYrbbxHBqWbBVXJFpx7BwbOZQzD3ZpFyLvRu8/6
VOx3Yyl1NGDxxnzpEKfSstHfL5dlrF7eNRvsGJfbyr1hBYvBt//X2URNs0iDLAx5
wIr1GRIphg2qFZ8ct1Ql4mvpSZgVZAjzqndHTYYtkzd13nULr0xB3tCS8306OFxj
DCXj1zeXbPRfjzw9WLFv2+Z0iUrzl1M4gqk4fsMNkrIcO8acRdV33d1IAZKVV2Am
ZHU8Q0yn+UIUbF1SU+0AL0BuBGtt4OZa9WfdbhlhaRsOvXFgsp1GfDsRqycwg5tJ
2FHtU38u08yQoHZ+wXupmn+r8zeaiGj3n68uo0kUCKuwhpxgPcTFKUSca1NW6wAJ
MiCcrT+N1HrMGkmsZKJ7hDFiUaWgnukbRCFX91UcHmTzEYS1wmUDLK7QcNPm9kXq
1TQ1/CHOGm1MrvPyyuQLjrTZUH4MW2IELOddA6dp+biGxl19N5yhtpAB6Qm7/dz/
nPfkbCz6y8XpRn7l5uNHY7nZ89GlmTAnDxZomEOHPyuBqhucgnrgfXbbnwLr54Po
bJdNtrRhJUcgwHiHEArDE/S2PpfoVCxbJp4hTtpycR4wyMjc1+xBzyz0fGrylFB+
+pleM126Y0216zHqkFyyY1ukLQyp4updaYUmBm6Fp9ERYHCOfWCcdZDdmHBmwcq6
akn3lbZ7StFIavCDV8AuBrHNYfgfzZgvcgr0LNhjXD7ZgfjLBBUStvnx6+r26c1P
I4H+sySNhVkK4lfmGaFoaT2LHWkzWztS5CNGbzqtR7Jm8B/XLL9KgQ5YqMDKsRiv
o1U0waHNLwpBhyO75JWJS+m0f52VkPeF2oszSWlxfBSv3I7spWlwt8ZV45LCnFJY
nhN/yKCyjsw4isTEA2mnXEC+RB2IVvkJKfstzvmVCK8Hy4F5kfyHRcmZXXll5/a6
UPIIbd9kNYa4fyaKKypsdc45jSGnszyp6U5osxyyb2llvXGHhL6LrECpK5HegvuT
z2VWFWGTLzECMdz1mHQ2lq+OMLmh4rl2998mrOrhKENtjzPXFrEdI9KmTP+OTAqO
a8osSUf84Q1a4IUWUPi6vzaLOEileEapfsqa1rvd7QkpGpLwujdvDwLQXH70oUs2
Evyp2ohZQHDQACdjyX5eAsiHQ2eJsFs1tbobTe2cFZifofyj42Sjiaj1jsXFFMsX
x8elVgULFU/aU10S5MWmKdxJzAWF4CMslBKCk93K/ZzTqyXdGtjzZB2YBJcZqQ5J
TMu7p1yCoxtwYrW15uTPBDVYjd5huU5KIcHnAPJU5ewNZEK9IhrdTWQe3FRic9ui
Q/RqaC19CzSUXXIpJ/7ngKk5y5pFa+f6FXMFuH2IpuIgfOMtlz/uZKwkrzk+Zhiy
3g8+cS6vz+tZ7YDRFkgxJTNnV3bILfoS2rdV1ByZ2EKQlOzJQ3x8eGJ8pXTGrUR3
AjGAobosfyOWTP28whzWUTG4Mty2bSBcz8zoRZVNTUzViVgBWU2nKppOYRSetYlr
Nj+faOOHOLN6ywdD1CCLzkpMvgFrrUxsfDOQulm1XN8QmjZqHsXFWy/QEtwUXU9j
PIRd3NDskrDfQu0jrTZKHHAoUgW6KW/dmP2QRUvnTgXVzWAM7tVZPXOVDDB9JWzU
62akFjWGGLzM9G0kw2R1oxxTxQNmXwFiF1i1yGbnlRPkRQahmm48uJjzc0kyi+14
flXtPo3G/EEAFW7rVSfbZDfAFwKHhdB16VYUkHesLOv0alXQ557Lmuf22shqRb0v
BQ5OHrsXWntIKCHXt3JNvlAQTlnYyscJvSjz8SJxAVBOmDjfFsNrzBNRo94DfKpY
NVbzjp6WecHG4+QqSFEaeC0FVoycdh7VJxHYaivsLH1PKGqLwwdFv+5Hb9lp6AN8
JtJ1M+b+iZGVduXCfyDdyUaIlyweQcsKntO+ha5wARhjATvetQb1R9m20weu5qQR
s0RfM8LsrQXun/3bqdvGcOLqQ1MaeYGgWh4Ygn3yBxgXUCAPXB+D8rAY7XRCOlRU
7sWALZcsNWmoqDoB6IkfVEWvRgMI8hIGInnsY4avEs7Fy0Q1OubKVwWX/sJ1atIv
kZaCrfeYrNeGxTtS4G7SQOs301IRyfa8L8hM2zHkHk6/RQyMqL9ni6SO7LL683hz
k+T05DZEHwVd4o6r+RS0HFv4LFt36XK8QMTuSSzSArz2Bnl9d9Pvik/cJKpOeIuY
nI9pKpHM19jLMJIHrBo4y7A1XYnMKZuufG2NRTSBR4tKVnB8JdRpwiO0sql1GaTq
DCTdMAfKOh3MSMrSG09PFMarHyxxDHXVyOHOVinO/FpwmL7vL0n28bxNcQa8ujYk
6BZCxP2O7qHZbNJzwd+g9JTt2RrcnVaPGkNbcWsYSAN5AL53QMPNLLKi1J2Be1dm
NRNI/5Z7kcD1vPzDcNdJcZV6bDuc+jM5KbvlfMrNihFDZlEQS0Zbt+AMCPschh59
1liSkki7hOBWneKiNyIffxVs/b7TsfmNYXHG17yPSq3055wIWyD3rt9FFegwyUhD
KoCtJRcDn/22IXSko5i7nZqXbo6h6XcKpjPtNhUKcJ33dPEW/2S6HyuGBypT7J2t
RIrIeuPB8s2oCmbBUeG59BXLemvCvlk2CWv5kacgHk+0bHGQyKGrzav3ausjIUuC
vnryWL3vgI5oXBVMkasWWDGXCDOcmdSSmHdeB9xIW6LGQy7HgY8+OyV1xTqbjcsA
ske2jkOii1+Obwa/vL+hcEFmgijdBF1olhn1EqSMh8RP0bvfKnuWD/ITw4II/Aea
kwwg9IoKp10AqZePMDuljI7hk8VJeZwbd6Y9uqyZ5JbB4aS2AErqIrNmy+7JC3k3
nRO9r7SzF/yT747emStQnmT0wSlbZDirmXlmbkiJvpbdQ5u1dWWSPdkYtfyVhUbu
s/MEZIUaiPT2tuGUtDeF914Lebrn+7aAppqzJRCNP4G/WBE6qTY5GGhzMJ94oAaL
Bk0/EeKdw3VbW6XGkGXhFdr/QE8Dyt/IhMfwKX5TTQCCXaCfpYZ8gRrNj1Z0jc3K
UiEJDlW0d6WZ7skGrx7d8bMmX2lTnkgbFPmmWt98LrOJPwOwOdn4Qy2KZPTTJh+e
OYpfG3SxkMtgt+sIrNeuBDsKe5JACEMimqhrhLOq7MvTUvT4c0g8esdYe2yx0GDV
TBkjtuFTz9w8W3cXYfHdhr8+qYMKJ78g1RXcfFvkb7errngwSRo4V5jOn9vVoWBb
Qb1HDvFdfqURbcspwIqq2ZxEbejvwkaoP/l+FuXYiXlzSmUHZ+sfjopjLBYCNXte
hMQl1dq9h68+yM3NovFwK854P3gTDxKAbVrZKONVarF99LgBcur32SDqQB3B6SMa
vSQHRC8ALb2b9nVZCUL5Ge8D9QWElv2THWJSeS3/J74qSUS0owaOP87JM4eQ/l3N
xHlTYrNIvHtC+V0t4xDkCYBYrP1ess0YnT7lpQ3kXo3uNOEVYqLjI7KbyI5w/063
QPvUeQLQTW7AEMHWD6bcKl+Hx8EKlUF5VBTbstAS59VXFMY64CNsBn6iwNnKn2qc
BkPYus4i7fGfXK/7968vpdCj7UXpRHz48iYEo7fvHZtH+19xJ4KM4F05tZieHQSM
mv3K/WM7nCXNvIy9unsC5M2TNR+sTEeGJIwPqBhJWRBe2Md7zOmQLiuJq4LD0sd0
mEgVtLBX3ZmYkHbHM/HHt0e4XU/w5LZ/M+Iix8PUolHfAOL3sv+DuHTeMj9GOH6A
fz5EftTRAzUtaR44r1/ic8RZ4secC5qfEKLLQzbFuFAtAHGggCHGjAUZiyq/1DXT
oRODOtaQLOe1dkRTExnL0bNCHaSEhgb9IcW+ZlnUUSDnu6RGkH8RTTEMKQ4K/VCi
UOdjkU37IiWnIqVF8OsxLqgxy5GKLs9ugyYxEdeiA7wY6uComHDbkm76GIZR8gZS
3wCP+Q25AckFst0pg8vFRKw+PD+d/D93magp04oKd+Vuo5o/olL43G4LSdUPjFGy
lJiPlP8MA9osJkOn/KnLNIlHpS3OSmlm8df3xGGQ3LGxxIn0B1g2RtNanu9inv1u
KZoOsed8eKvJlD30RWSasupDF1U+1TQu/BABvKReLQA0VJyWhP9wgx/21vkSZSs5
RxxHH86SPVXH2AhNIqan8sxyQgq+iV/TSdag+N4jozE1yyM6wZ94uUGVJwjeddU5
MHPRkX9l9U1BewLYDv43crfakc5R2f2baBV3+IwURUdVVGhe3beSKZ5uZMbH9E6D
2He8e1CUiDbb/adrz1to1uIPHJI+pzoTYE5VoLj7QRdW7bwOEzroAhkQ8apWA/sm
r51Y+Or7rxzsZeR2FaJaZUUuB5FqLXRy38Hyn03WylA18hCLeBDCo1Q7tqJ2NrT8
9VYPATrHqqwwHxPgDYV0n9KI6z7T4P0ZCoWDGUn9NmnqjuOFqLrOgE3c72omj6Sq
ORaZerL0lWsJV8AdgaYR9TG83CZn9cWOzLbNm86PgTjdjy3bcL7tOCkk/4OQHKo9
x6bVdQEcFx6y9Wkq7WWXkGHbNg2e7IA78sG+VcznxNfQkqBMtEa7jRTZbMPOYn27
DYztzg5M2MHuF1N5rcF1DPKXxTWUoExVfuuGmwkyEGKWYA69zTXIJR/6h4nQP4hg
LkF4l6F//H+YdOUb7hA1xtIkaJ281LtmCLP44sWg7tXRsh+i4lmsV9Z+H4t/s3Kt
sJq3O1P4BH49g5h4plwTJh5mxlPyNZYnoM14P8Zlibo59i2tn4LpynKVObrhWSF0
jMRY5wYcW2IDjXW8j+w9eDadx9UwX9QfRO7Uhcb/oDYWLen/oG+bCTZlGruHgdiR
ioYgy1D38KKEl4ZZf28qQFP9ZxvkPWCC5uMcyA8p7BBvwmvQkGouVbrKjboK+kyI
fTtGsgJkksKrtr1BdIbfpXtH95+QWTfTQ1YacPyQv1TqtPBADFCRjNHXxDZJdYvc
mlB0O93cY0HYsq/ljZWUz6Kr/XnGdc+IYSsgA1oOYZ067nnpm2xRcBSXi8+MjqvZ
tTxoralls+AxaPNGU6FRod6iEd7rGTq3w6XSFJ1Q6BCJvUAO3bPjikRkVownX7a+
P4UPOoFYjiHllrS+e7aCiFdCs0vgzmaBNOXzJWEJGqa4sNEpSPGJm2QPe4UEQP6b
bBt9j+RzJ0VZCicTZe90XDtA1XxQ41169SKc6Ri4Po6J9ZGyD9mz6nJz9DErlLf0
D4So2l7ekVY/4Arh5vA2xrH9p3JA6Lr521HEgJDT487v5K0axqbIowjXQAwhWqc9
i52sQO5k62GlnY9jIKJcON7Q+i1mbmaXSu37OyUY5Ze+u1YEnwv58xmmDeqoRm0v
EHXqGIwgXU1N/FVKn5dW1lDQ+vnZ4/8nOTD1bmDZcf0tb+AlidLvBKosaPsLzxXr
NRBCLnuuPkrN4dfYVHM3dQ0a7l8KOWUSOVIwa8ril+fSb00FVLZXHHtlIvlYOb3f
iKltdzTVSsEF/XI2F9DdPRIB9kSADM7In3tpjUHTvaELypwANnowkxA+hGqwMclh
`pragma protect end_protected
