// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:33 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Cj5bk65y1pAZ1uz5XLkSZukogElamOwAy1A9SN8fNv4PBqo2yofQfmin0naJfvBo
sj95mfsMRBTRn7fpPGB2OlH1DUgWAL9c8bTlrVDDft3ITa519t0Eir2ca0FDAnhF
A4TbWQGkCTYz27mZol/6nQ7opuDPYdIJLpxOTW7NEes=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4416)
Q0oYlMHkwvz0NMip4cM5byH/5qYWblAeExvMWPh4Yg2DhL5vwN+QoDskH9WfE01v
bCI6nwQn8A9zNLrhwRCj8ZSA5zT4gAkL1RrS9qcupI5jzDHw8xpaVntcIA8CiZiR
SVT+4kq/GVEfEtOjalZRKG5uRdHFgC4NkMD8zTorw9LvzQ64ZhTk8E5gva3Tlc9s
qQoNcycXCy2r0I1bpgyru+KG7sawr5qCix/WfPfvYAy+cpFwkH9njeLApVhl2xID
VcijAG+Bb796BeD6ltytoDiM3nYxJI75IfrwozJtL4K/H2MmB6Pf9/y0eL6h1bnO
W+XS9VyE9dGNq6Hw4AT9/8DMqZG264ygfRTa7p1lLZJDWBSwOWui8aXmYZBwQfBc
znjfaqJ52D8k5woP1VuNzdtkrX+1H2Xft/241pYSFbN9NpenOxmLh0GAmiP+UpRh
18sAT6pVU69iUA3VEw3BF+DfbcVc4qlDIVDo0VdlF7TqyFuJlKixYFh5nDUX405i
0vIdjx5nTMksKSzHM08HENz60T4qlG804D1kO+e4u0PQJKoJ1ksRjF/1IntDWiVI
8vw58kfV3po/nhARfGGDpojbE+9lj0AUALluxQraQg2xLkj/Gi9tyoJD7AWWMB6a
xsdqQqj5LRHZsDcNBt3hZ/aEGYxsXYhCmYoGE4Gq3Qr5gXBi3m7Kh4focLbTaeZJ
whywZJcJsjgzEqtDdfRWWEjSf3l7brZdaZ/u0e4F+0y7W1qkX/N9E3qb0fK6mDu/
4238OWeKhBRj7Rom3/8s9wAYSbwrmp/+aq33tEWX4NUVmKYOH12hjA14FX2Z7fb5
dbwTcn0HkqfPhi4lPIo3r6vzKQQCgL8W8ZJS7iTrPxAF2Muu7NRJ0tkgdx5YUVVX
l1JpHNb1A/bZ5mU7hYqWKxwc+amgXe9LcTHHhsaPgMrWENpkfAIw99xBWFJE81Mq
mKcx9xJPx3ooWbkYxNgqGVIXJZbAziEB9U/qKEWhm7nc0ubkR+QawYe7oouWhSM4
0U6Fr9atXgk2VMhKtHN6J0eo4zEdLRQZSVd11IB7VuCj7+NhPozix7zNXPrXcMIY
e+2oa0Q4yfeuQrpcOocBWRApToPhtzO5ktN3kWXxgvd92qVVnBCAxfYyQmfUE/L/
HRnXzu8zimN2opphL/GvUvuSctuXejJvtdtDdXp3nUl7Ug5mNcu0Q1YoVhfAvKQh
ctxHPVgfADrPbiaK2qhyalw7dd5AZWaRN+/THY+sWyj/Lrv5KcxlzuhhfVCGqKqM
YPiKEQeMoMxnv+e3qIqNO9kyHMN/JM9oW1LT4y0ea74JHQCGYCRVb/Uh60ZZ8C9I
pC+hVq1k39TKPQgJqrCLWwGXCEpUTHk9aMkXwweOtPapf5kdeJwFy+iNrWto2kBV
GG6f6Z/Oz9EDH/QIykLsxLuvxeJajRY+IHGlwc504l+f5/+aI+VTICQuK6LkUmjD
7mtXPYRiABDAge+Obi5hxu3gr6AGAV92dhIbR1UBHp9MGoYX0st1Ev5xh6gnmBdQ
vHhCzVPWkP5nMTrZzKFSfHp8M2ZY/bdwmecCL8LPTqqEY8pY6XPLyqa/9HU4LzyJ
pb8FEPyRDWLH3cqqToHOfvs3ipdLO4NC0draDOogvFSgOlEiOXu55K1VzGnDjmbx
9lGl5LGC7Vlw3R/mrQYXxDIoWdAXVTdSSifi14iJi58GxbxBw14taT04XQILBZzY
2Ug1D2CnfQhl0aIwE7vkQtTCl8SSNV1lsgyrN9ypiNHWHS+POe82E+JFXahyT2mF
Z8yU0sMVkfH7fzXQFvCv8B6c1Fkg4xMkuJA6cie38l1GnW32gf1GGoYP5u6A0wcX
eSPOg8tPF9XvhzqOnu/KZ9mETzMwgWo4pE6dYL1WPsd0o5QrjRDmRjIz1HRjonTM
aOdMBBSF+DCS//4gEUtYdWZTMjpNd4cGmcPUJ53MKztqPAmZSUWDjQIShYvH/ggf
jo14cPbpDLOKehXbtxYa/JpKUgzlXBzCsWh5STkqp2XJV+iLD7d3S0HHSYA0c1pg
rcVVuTb/3xoXQ6F0jCZTUyZAzL8oJh2e9XsGenwzfhfZZZhddGoOkmZZgmmqRqM6
aXU8AKOZtTC4B2yAHdbgtJBPt+MmG7jkp8+YbqxEsmURvst7wizhdXi7p1km4L4Y
c8nu0EieuKKvxt51tknd85LkmQeV4D2z7ULh/vM10ukWTVLTGL7zPN0bAMlVS8fJ
BUxs3ue14FNI2nyIoThERwzp1hie40WHKwPn3HoPahbYR612WwI5YgnVSFnMUJ80
LmyYrOHYMtkj+jU85Un5rJ+2uWzhvNEIpGsgePJKIVimt9uk3fsNlEh3F3z6ZQT1
qtw/+67ncYPSTi9r9t4gW7SEYi/bAuFduFj/IBWWYFPeQB7qVdUyamEgYDzG+iio
1Rc2v6xGXFulwU6TpTB1X8FlauMlArCFruFL3atXOGBYuaOmqYXwJqPia4YiiF3S
h2BdHau3XruwpWIwEsIhgTdKLwu60Up3WciUWGOvjfewfOmKFlNKKLHiP/vX6hTe
j25SuKM9sI7l3UGCutEJUslb4K5nGR+2OSsK7TN45m7xqNO4N9UnEmvY56VOpS7+
2kEHoJCgfBnh8K7HDKRYCWvZmnyweuJ4GRint20TUPlfyWvc4Uts8zv8+JsL8VYn
YRIswgBQbkplkifUUYcrP0xMIGqbpWvDcMCi2PNYZD0DY9AjuenJPJWGnT1UkUYw
osouNbyztXhfHI2cAmUYBo4wgy6OXFHS68DHbLf2n6YAQyu99DbV3vH9jUarK7nq
gO6atWls9fUiARU5dEtxNWsoAXP56IK+gYTQOCiEosfCkMJAw8vely28VxzkJHCB
FFzlijFWwaH2JYGx53T0CBZ0kUYU2R26rzkCQML2PFTEvqkhBj8m5XxiUTJET7dW
JMeK1uCLKjN/+RANwpXhy76gdVlCxrSRkTklsqx9qBaImhxn4mVeola8EGUuh9CP
q7c98XUSBNZPQpfiUyxSySVWmo+l+4Oe5gsLLsN7+ITRQ/0CJwlcXaM8pJvdbdky
OiBxeOEeOvnS/nBpgSY1sT5upjizSHLlQa6ZqHMKKfPsBNS/zmEa/IrVOVWOqXb1
bjWOh2CDrKeBdAvwrIhNHzhEfszVRx+ffYi/42h524AmoDeebeA51SA0TZzvtc1K
ABO4XpbJflIQjIAZID3xRbm5ohLRksSScxZMO0xRc+bzhf7A1h8N/T1r5/FjG6kX
9ooJg1nA/uE1CXTxzUiV0BnJNTIedHIjSPY37exb1i4Gqjy0ktkI1WqDoT7D7LNi
ko2oUHhy9KzEqtAlrc36ZXZ1GiW+8a1n17zMNTQ7CTJAVU7+iWq0XAzmD6P3YonL
Lu0oH4Ed4tZ6b2t1Ep+p/Rit/z++A7diJCc4EgF4l0SyZ/H030FXl8fodR9tws55
KptkxVKCXPS21I1w5W/kErzyf9m7EA1HD9B7hx7ByQON2P5Gejp7Bpl8u4TC1j9p
Wc2ZP5Q0nnJaJkTJ99Pi2a1/FxA/gxJx7drC8rTwGbp/stMw6+VGVoORhJoFeysz
i0+lOQn4fc5r+2cOQMwpJIdMewzlsJ1nSDaxfOpnT9vFScxYdzHRiGpUtht8V8au
Pn15nxfSQ1KGGQlGEXOotQJOA154PgJyxLutt2F29fm0gJuvA/Luj31A9g9g6pOQ
mbTOqRpKQa318L4Qqa2/qRVD5eaoJDabe7FXksSF7bQa18T23idOoaLJHriBkmzA
ppcqeSHoMEPvTONySfND8pwTOyRsW+r9yAezzzsk0cbXIr9Fp9BBoQdezlo1J2Z5
RL/S4XAuuE/PMfYxOOX+s2buFiZ5LsKbeAjzl2A2k/98i2ILhOaN4BFtiEKZFQua
RRUOudnMcuBtC0owMszwSF/8tcPRPu53Ci/NyGIoRjSrmAo1fYp3XSrW/b9FrCJK
X1J9008AaBYhPd2wGGcP9rvN6jmbJd002iCGdxjo9UnSgkADdsUnPlLYKs3+CmMf
02fgXLqMQ0UlCoJATr0Sn1j70fZTakGwBRUOPlnqvdYcpMc+WLjT+Pedfqz5872X
s8BGsgwRAuu6dP7DVGIQ3YjRyWvIqMUW14Kny7AgopnM1zSN34CX/AOt1IJIIpya
0VoXgsgdcCG8sqZhXV2I0RlZ92efaN+XWPYUKNIA+nZ8Gxl5cot3LXU2jvlWrbQv
ZrCnk8MhD802EqajCEaWuJ5CMOQwelbw27h72mKM2f0a9CyjkkzCfQW2Po/4MKGm
xy+iOhLrDlCZviDtBXDoM6ybYvaukeEieah9PT2WbsOLpBo4YsSQYvM++cNRXx5z
U2WmBfO2b4iIuKTlqtbBLW2clwtK3fcioM4VfDleL8acQ0Qmzrzi2AhmlDCdPyPV
6qv1ETzBAv3w2NMfbelgxbhmQA4UEkqRbpIdo2eLvVuxbVcYH09r2trLX8Y0oCm2
jCMuSuYtgmVdR7QsTRvJo0j6MSWA2v+9SlqdWUvTOTTfT/weZPBq7oqoRxOAHunT
+m+H4PDFty7ot3jgj2DKe9UA92PKIUhJLGsQmyzcmTCz4S19nXX/a92+gi/TnjG5
mR3y2EZuBMBiJDGI7uJ9XmO6YEwFyh3yAyW8jQXLkl1WjJ3qfH+2cZ/8dYZ2JbTe
yfvzRXXoY5GXeCbBDzFPt1g7ksfscWkUIo3fbV4q09BbIGTn29liHxtmKaQqfz/8
eiqkerpO+qCDkHTFFLy8sO19+39ehMnn9KKTxlxit13QPuCNfOQ7PUxoff8TA7j8
CfV7jYwjymAVghHQe8BK4rbc1UtQMp/3qKSkanipsUxD5nOLaIxwHgx0FPGGNUT2
Mrp1Ywx/H8oNPmaNqildTKdX4L7ah7xG75WijBMZFBrcszy1drqs/idJisq/k5yr
jSUeRsSx8Yz5IrYeNEEJh11unqRIENrFiJ/xKkL3RUP6x3FWfvx/p81wDG833Rp/
9Z6L/kD0opk8+VEJSCDBzEidFJWmNc9AYBnQUndswTm0RFhkhZvA5q+Pv4GD2wxI
7XZnzrfns8gNX3+x1J1oN3FA4zOKydcOG3RkeWyR9cMMm8pAQfqYqWrQHcqXn9hf
VADvBaoM9ndbYYgtcsb3PquuCgVSYIhA2hSYjVa5LHvIv6Lvtf0xbKZNIgGu5Xgu
3bwL23KjIeW9HLnSwjLGU6jXgv8tD4hERnKWaPFf9vOCkm+IpRKap7ElMlwmTNGO
PsNtXhxvQ5DgtvfDzUAAEN33tCYk6sd7we+BeABY2rzHZUq2HK5pvRZjbUtXX/h6
pzVefoYDcRk1t0L5RZo3w+W273e9WuL/Vb+Lc4BoXGFD7vLUmLHIyNjgvG6+cj3N
jQ9GbwYriioX8IJr7T58VNkhVY4aH/JusW5gBEciygi9m4ke/vNqqs/vnPzTQqb0
YKO3xgc56nNOlAxCplnjlvlfAvwiHFEVWXf4OjTxOTcIwyib0HLbJfrBP1e36nkZ
RPdykayuR78e9eHGrVCSOORzHk0QiPeEfd0VpnpcBtuCpUzLAsJPlNpDIicBqwL+
WLBwkcOyPUW1ASHy1geb15c8pctwz77DCpyOhBHpqMobYS/o+HfnEUISELUdyO56
oOHF1kXE7Vn0k3r94SdfQmtMZUIcj+F6q7UWhfQ7pQ434roH9RNvaoZZwT/L0HoS
L1lk+NP3+/ColKq0vlnyy1TORun2oa61HxgZgWVnjh5sKoTc+zg+8dedcSao62Yg
FEbcUlkVkU9QAVsEZSYpS4c9unVpmJrSBJFxdtO1hUs7pTIofrwH+lwWzFk8uGwG
DFAJmuBw8LjAiuDwgC5sJJ8aXdh4NBQeyAqEd01Nd4pxH1vlgOlAqm7fqv0vKjcp
`pragma protect end_protected
