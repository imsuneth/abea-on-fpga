// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:43 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K4uH/OuHWKsHHXlCmJOfpD9VlqAbPyvTGrogFku5eZPSkcURM+9yU9DvoJiI9Ywx
x7RJFFwDTMZVQUYTvuh2PbJZZkthPzQ0m9CycggJHWqELlUxerr19Hjuxy1u3pAa
OMQJ1dKF27qxGsCujm/QCUgD8A211kxhagDxr3IY5Gs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
FaUTYe/5IMXV9JIjmMoY5ehjrT1TpVgt4lMDlgFHk4G9UBA/9g8MSa9+HSrsqy0X
F3M6Y1JvWKEg7COnTsnnhy4CzvULOta55JJofuR6AF4IlKI3TNoPXSEsJWqOjujr
JBXRE0NqPC1Xa8oAPF5ORM/9pqWAaO+1heSRwWKvj52FFkwchpS3pjPxxRG9MWFv
TGl+7pLuM7TkTdABvhMWpu74jd8hnGbNwfB0evIi34NtnOntZInttMSw1GKrJ7Ey
fNfF9z2kow77QQJnInE/uxNi9Yo+6neXVwEOxF1LyDy30XgFBHXD3pXFP7yRTSLb
afWd3/y4Htu1vVohvRNWGUe9izvY6OAm30P7ZOJhWhbOhpthJSPsnIvj1ne/MFoP
ci/DiFGkR1LJidsz5c054rE+HIckrUISX+MtJj+sK69ZenleSAf8AYFwyRQeWd91
jqubyhzJZmqe2QpntzBBU/mpGBTXfmazRk0uPC6T1UHiFmrzQjvkUrmdHryvGshK
W28idfpzdBOgHXIh7k/H+NPYxjjbPUGaCdLhMmhxAb0uBMwSqOUPpUePOOdV8QUu
Y73GTTmrVC1aTUvkXN7YO8wxfXKn6r1ZucVUAUmfy8H9Px0helG/9vgK5n3ehzfH
L+BqNWunn81qCRoZCy1Gq5Kr3PD0FLgx2zDD/ncnwLaisbigm2toqhZexyRpX69t
n+YAFIXNKLTTTG7n6qWvguUqAQLfV6ubbQELSfqXMPBFMKfANf7F2fuUOQoL4qEJ
VcXCAyiX6AkmNdO/pXTPR8ye1548tClRv5+spKSamo3vQDnxU3NFprNR8RQpKNhP
hZeXSSeEzbcczBCNIJk43dHoycurm/4SX6LzYhmTglM1bmgDBi2DZmn88+JEuFuH
INhhXmgLu4seLuXNopI08BD0tZv2mqOzxOJY5CFKvNCW030rj26ZfqAx/TrhNR/E
j5pJZ6/Ly3ZpyWFXT3mf0DlinViiUvE4e5UpgHhSiEsl361IASxUYEbjx7UELLjz
ID9xk1wR91SNs8x0WCFKD0jlSOycY4QuJ692M34AaZKy4jVt6xcc3xbpMsIS2XGP
fcfWhuBaqJjtneK0/lLfCCXU9OGq/LwDPvrj960/ESJcv3niDqrZ2GZ2jMV/rxtj
ggTubNEJfm13zIXXmG/XZUdP7Ew0cGG4lMu3BIN7wEv/RwlYuMR9GUASVT+1o/wF
bJc8VMeNMJEGxEaW3xRcp0deTQDVwZn+C29f3rvPgPcET5bVDtUic0gCu6SsBnBX
GoxrWuUlim2i23Z8SKvtc2FJz+9MXkJjZ7QeV9Tw+BSmacCEWaykQcvzHyFnVnkU
eYwr2pmJSEiysqNzkiS4M3bUOx4iy8sK9PbsTFm+EBP1kKHT8Bja8Ncs/twxlia3
x7H1j9W5eSbEh7WD9plZmFMuxHyHEdJbqXZm/QbRskzdOQabMSSHxDjBynl/rqhg
W9CwzVpuAPBcN4oHqp0Wr2IeMW2yP9DZtqgWftTp/c7tiRKUZ1zBKcITxfuTT5Bd
2lB0q/EKN/WW+8UiePFqEnsly8RtR+SmpJDC2YCqEJFnVYNdsz+j4tIEGLx+2/uv
rwHpN9+6UCODvVDWGvAsv3egtipu/jO4Gtvl6AJzeJwy/vwNEh7c0pkYN7J+BgGX
Sv8Ap5danGpD7/ScFKrEuSecOBMp/N0PKIrVQGvir2rCm2qNQ3Xpcf0ytYvDtY15
1b+sYoCy/4LRfSoTrXg1TbGDYaLdlnOr6oiPfvLo4OWqZmAwm85tpgig9cA3gifj
oo0T9iDxGici/2AVD4BYWGwlVhWT/y5IXmCsWUoNknVOYtCZcUTfBZ1sIvf4UBcu
djKyn97/FJJ6dHsH0XMzl5Tz3IYK8vjoAubPBmkyVimr6NFaY6DKyLJ8iKsfN3L/
ZtIfizqBYAN6x893fi51PCsHoMVG6EWpTvAj/wC0/psK5tOCWjNUrvaA8SdqZ+qP
VaclMoxl86FjJEv7hWdtkESrNO8E7puNy5sGOFfOOYBOoR6RXK6n6izijKNO+5ma
AkqrAO+kH7bBxP8y8xhGPG8/aecQNIKK4ci0kHaKGD9c04Op3pp0J+cxLd/LmWqc
Opr/W3NhFiDbT9xmwwiAywKEdzk3debJhsUQL+Dq9jia5K0dH0tgcsPxAeT6cbGb
3QrNaYMJfTNWWulLCH/phpP6dHQo6pyWDZK3ssO+698cbFFl+CgVKTftQahDcOnS
U4KXIXoyWkCiCnq4aeNP3p2tzjL4ZgX676hKOVmcgisTDwlsdvXUdpCixkxIrFGM
NydtSgDsYTe5UAEMZ6SfZ8hegNIn3HSXXM6of3NGTdNpMSSmVFhA+IK7DN2OLFMf
MzOW1xY0ZXmHCht+Jtrci81I7av8Ilt+MMwNaB4bN/A6TMG2FCBoDE5x/dAsIZqa
p9KxCvQbOfVDbd3pHTYd8YNtrqDvUI0C3SpiNYK173d5WqenZ5fz5jrGt3dE2Bpn
qvLLuJYEHHWTHu42vDakpUBxOxLgXhWzGuxDwXiypKH8d41yQUOwl6IxYnhSp4dc
1h5YpDRqBjSvbph0miP9Mh0UpEiEKSUat+j5MkAXIsW7hJYpDhJuah/Rxp8zI+Xl
ifL9gFiqeg/g/16dfLQQWDYgXqE+L0HINc8kk4+PZ+3cENyvXxOXj2SrP3IlTSeQ
dYFSVZNi9yyyh4oJMOjF8Qn3EdclEqjoKO5Tb0kF510HDaxnRIk+GyhPnvkwWlZ1
2RG45lFQsWUa9N+SRfaX2RoGEn42NDsVUW4WStL1I1WmgvpeQPGKfyLYKA9OfTOI
SowWZwGPBkNEhPBq2iFgVdJkDb6Qjjl1LgQuu+GbBZqDCZruDINlju/UooXM0r00
Oe1/D3SXRs7/hxnymOjC3GKeF1Lp2EfCbGHUdgn9NZZvCRLVDA/TVIeh+pQbAEOM
6CV4UWAGvGOl2oHU78A2dfpLIn3gCB4C/PZTsDC0VhHN1TdGP/mhzmZv5f60Bogy
sps1qnhaMTpTXCJyYAYxsCK36Wl9c5mxovLza95sDsTWwLSuVp6MP6yXszJHYIOu
IC8Xn5RNRuR3AonoMy6Fxm57CBv2c6UACjlMhEl5wmEwa2PWMtJrLK+chx4kf22z
PHEkb/KPb+hEiFiQ0dlJDTPh2AjkK13vV44/tJnAwzuts1OzZBrKasyzqcTs0Isc
qLlvLh07Vekv6Zs5PpxJ0TA0AS8dcVXDsiQ1NkKf2fwof+2Oh3UeHnD2NPcwoUlW
cCOD/w8ic5deR8rVo8+TXYr/SSsIvvbQng16Nz3WuYzCO8FA8j45ahlmtMX6whFU
0SNhi+Ibqm1MAYRA5DwfrZ/zNWo7CyUUonIjB2CYoqDybLxVNCqBEjjK8vzE0Sw+
G7MNopk9UDNAjkEdyqMCpH/1DfyjXxTUijPOxYR4B0GEbkRsb7dlludtJwpi7UsU
o3oj7C77KPVJTMwMRik5gZb1VT3gt5b7lHgaicZeiOC6kBY+Qafgfr6uh6G65+op
AT2CVobmL0z7tNHxkiJKMXtlMcc3JeZQbpsKO4f2aioBRitdKz5Cc+Z3Sdnufkvp
wcYhKNMSsGaFYKqIsqGjxwkKE8ugF3brDEYUQoosvjONEog6ygJFlM8y5EyEz9DI
8Cs4/4CwOILDH+exkH7QauLXcO9ee3KrX/pYMfVYGveLOvMH2xbo+sCc3i4diava
tiH2SYZRNrraukiQcKeELxQWwz0v0EVd8CnTHz66XWy/CqvQ9b1IjH1UuhZeoS+s
J6VZGVbV0dysy4zotOx6R8UcM7hO+Lktxb3gHR0Uvg2rJGFglNCJZGdYdYsizcKP
3fYHehwOnL14fjhi5QJDX4nnf15LP++XOfDByohAMV1VCuTM6Wheb8iB6aNLxsAX
iKGDKkKhUI61reg3CrwJYUd8ld8LXzP+fRMowQ5MZ/Ej5pbB6HWSMDWXs+Blfb13
dEtws9cBWEzkJLdmTaUHzYhFXmQUxwki29stgsxTHfITpZr7khp+l1KsoHnXqMu9
jxCFSwplUh+tNqs9Fcp/5w==
`pragma protect end_protected
