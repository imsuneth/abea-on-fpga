// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:49 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QmSYooFYYycjTkKGj37nTxJq1OSkKideYSAtTS2BInwqtumQ9iTl8OJRhTVovuJS
1qbfNQLmRnwxcr8hZCnsIOBXcKx2fMRBQVj2hyD4dpCGpBlWN1bqKj6IHx3KW26s
OKYFyjuijJ81Yhs8BSHWQBoFOnf4QeMpOd7gkAs+Wvg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20160)
AtTlXZdF/2F808H2+xy/zsE6bbK/5obe+gwGe7W/OUKF5HyZxybi480+hdB2+Cg3
kVgVY8qBv1gx7TBhaw+iDz6Kc290vefH9FBXsmEAAR4r6097BX7yqo0/Wh31wFkE
b1tXgRUpKi5METmLAo9+Auw4cON6GQkQv2OOPHf+KjisFkUjHuVnHU5zfu5hoqVC
otPabAF72On0KRS38zggTuf+Zx86brBqP/Z8SFB5K7lU4OnLMJQsWseMzgi2IG2K
o7LnbJwLg7UAADps6t5ZO4UvYXSLlIlSZl+EDkebRcXOnJwo/q/xGfBMzTm1mhNQ
vQ5i/CQhcXjExloHiV8t1RrjeZHDt4O7DwtHwkVHtfqQ+8VwhXm52JHznlMFPR6z
BiJ5fI4SAdjHwXW5tKOmey5U8+M0t8bQWG5QTYEPEtkhxuvAaeFyqs9xk+t4NsIs
ZFMH2LSqyVWGJAZDsGv2JbdFZYUYEwenOMCHzmc3n61OGQ2lMIHN+SM+Gtv0xg2P
rOHDhx9IhkRERbH3ptWNrocyAzkvuy65GedG8XBxzBGKddnJi1XuPhiTsz4dZ1mI
/sB2kA/WH4Uwprp4n60x3gxQGPYskYHYYCCpiR/wwOYZ/vc7Y6h1KnQzov5dK8HC
hgLL9GhXyMh5vhHQfTPK6t/voy8al9KnN6oM89ZgEKqcir8Igoyq6AZ1pqV3/x/b
AYjUZlsPwXpngmSKKnhzSvZFADIl2RYC0uLI+mtI1ecugwpeFL5GRBrLIc9RGHTy
na0tr1g44P0yVSypAe7IUYd+pNm4srQqIvWKUd3jbr6Qzxt3thzFRIM399V6z/MP
A/RwkgtIwKDC/5KYmPh6fNT0zBXXrAeh90RsktoRLdmCdk/d46TezES4FsQrCxPq
gQ19BKEnQPG6dAomEhwZTmBe4w7nRfJ05R2Ga0mUfAxH+B9eHnJfy/eQlLvPrPjW
3wOuWrpAKpi1/HS9ekJlJX9yzD+WRtAJ0R4e2dIOwCuTrP3o63rLv2wnrFTdj98R
Jigk74Ld3CQSc4mwv/ffRLz902g7+x7ajcA/22yTOtSu+TbanPZVZ+4k9a/FpH4+
epSxbw/1B7bxggeleDjpZlnlEZH/6f/bTDZaMQDdv0bpF2tb8ETeE7l0C0IuLeLM
32/gCif95xrMIJwxhrIdpWGJvdy6mQhMyEt96L7RAt7je5PcoZJAwEBfis+Yzopt
4ZvxXdweLzftn03RVnStmjMqD8HSv2o9wF/AhzQAVFxuZsm+h5lLOyZ+UzrUMv5n
5JNzCP8fxRDWpNcKoEVVx93U24UzHyzvBHFTrUL6n7sssfx8gjd10jarM59mTqAI
xL+DkdeZj3f32jz+wZyrfbhq4xAulSNa3EHJMVF853TknTiboIxddMAg2FIwECAF
W0pIGWNNErJjdb5/grE6ntL+55f35Ci50iRDiOWj1vxnEsHhw6GaEazoMuDyZsqO
U4WEwCJldUXE6dHBQ1YufA8SBmxxATjuzU04VB3716qwoL+ML/aRm193r19UwK/X
hvyZkhitcOw5rbmHuUsGtrQbV6mmBPDkVPGqPWcZBOnohSvlxLvKqxg3XYJ/2DmT
RHKC9N5KGTrPO4O/77N91fM3JOe/+6PHPMJCqWH/6CzEKRTFj4i6p281tBW4TwNq
GDEWxCFy89jf3t3uaJxOu8lqAVMKJA69jxNXbtzWAudDV4ehqWGnwG8JEO1jRaIh
x6jJ12vGtoOFfzny/9pBjNpSkho2q7gprIjfOMdFttqUfRLMuz5KIMqOBpAoit1K
QABSgc6G1PMcip+n3rM++L25aJ49PUDadDZOUcEfne3H3FxeD8McDWLbNGQRBPT1
dbp+iM35hlVlBZP4Fah+jbvRnZexEsN1gaw22rIB8t4c3PnnTs1UAO6RGza/rT0q
zti9RaGG1iH+6+4WF8V2E46OeyQYySJ0Oh8Cihq91JMeI1dB0A+3sw0+04Fn1fID
7DoiNmEApu+DtJpx9kilZgeWWk3h0wVw7esojqUYV4ToFOqC9YVgrZ/pqT1A50MO
4WL/0+bCiMIzMdfByjD5ghzz6jntay0yIUemTWHa7zYPuwe3LU3qpgIITc0l2aUi
3y3mzxwZU6gOxhlZcgVC+uDlWywqnLbZk5UN3OJxYGE7YoObuxPl2FsIEXaqmIFs
sb6/v06OlD8p4lutPX4heDd1cBy2ajuuo/HjT085vhKQ22tnpwMrPe8kWXJ6BnkG
hs5QbfDOYDNuQfg4SnxmdU5sLEc8+iXa3feqo/y6AX5mwEUbI9LMGXrGskhoqAya
kFLl4gORTnF++beYVq47SsHTA40hQco/M1f0+9YV4pGuUX7DzLP+R3JnG97p7FRZ
0orb15Va7vN4ndOr/yqhhyJhz49iIakca2nprsnTdJnIfzzmODLCUlEvh89nLkFr
ZQC/66m0esPgx0oTBLpvKBu5ZTdsUo0jQBRzkIcSWm3J5kJCwGOdO3Az6j7Isj4b
qgKy3UJlKfG8flQRcKphIabRQCmxJDmsBUVuhI30h6AC0JmLCX6XMo95znwHfCIw
1QTthfTHeuOtPfxHEhmKe6lGHTpJdoiVoPxFOMbos+v9Jhlz8cRXEcXd15zhR/Hc
1WjyG+CWpCniRUmWeZ77BgG0oQbk6VKCDt1TeoJXh5cfZvKidY7HVu4wllfwH7aT
mt0TowBjWGts47vcUSqWtvKjl7iVeFnwnyXOUGa2i/38O2RtIDsLSmKRbgQVIYR8
xe6DQX7wJL64CKtTOx24VOuC8xsko0+8pOoFTkvS/9db5ZzTs8bLdX0NUk0HR8RB
rtBrVenKoTO1Rq8bb4VNKIKDO7Rqa9dfHngCCRMqzx+Axu7ejfkENjky4zyNarmS
RzcUGNIOnyCks1j+ZqXPY0mdcU7AQ0KChPyZIQgQZjQiDge+YWiAJt6mGstKEhxf
pvLZ8ivt5mpOTDgN2sdP8eOOqBDR9AG12+EtoPd7hbbbBI3f8Mnq40evr6/AvapA
VkMLtJfW4LHCHncVFkXtuG6xu6zB4x28iLYpqmtAlAYvge8vEffad6Dm+hIvDjZi
uFBObET/mvqMdGP1cyNqSEZ79q3xJDx314cMAUj9Zo4E5NwE/3DCQwQFkbrGEj2o
1fj6oWafi3bKp27idCxfhk0EzHIcx8dGy6jhr4mTizQmnamezx7fzJvj8Papk1RE
Dc4ZcD2QuIht9sTprnSJYNRXxN5cMakXMUylq7l+I0u5vFxbH9yIVFysMWFVMk5v
tVk5Bxbmp7eBUphMtkNEAR+PAZOCOiybaHzhbkPV+mP2CiEL++tI2rQ0UgXWaeJY
2+yvTpCUivCNsizwoc93/DgkognsRLvskwJH9siOeD+hJd9dD89SoyM2CQdxZKTP
cKS09IFMzY6g2nzp/XeXePp50DDpEthVswm3rzB4z/CoUayUsmeqVAKj0xGnGNjv
C2JdYK1abeCb4mdlPx6BRp7TokbtF/4B8E/w0iZxxaA7lEc7KekJoA5fjZjjbb0i
PrV/PeabAHGYCz/7Nv640h4HXKMzOEgNw7HhVRIPEnV16sP+I+Z+q9vbuPXwOi1M
nwPkH/I52oXVvn+sPbW0A9MKXoQZq87QD3ASnJNHJqZTaPCESpSTLSefHsLKA1oo
98rzP4oZiRWNeA57bRPn67r8k4mcq8IPQcUji5FeqXKmnuOcsPPoJBZo2CAakKps
5UPhN+m2vFeX/qF48dzN1pGXAZFqwdORp5MzWIw3Re+V5gowL3ZhvppxFrVccdPr
97uFNiWTp02Ejn6pW3rQZJ5SFr7hCoEj5MdEAcQVrGeEPa/gSvrO2E0YEU1bW67k
TG09ccx7RAA1md9G5Y362vFZhK57s5fn3nCzi4UQ6eTyOC5wzoO70TyDTdZOxili
tIe8H2Kei0xN/h4mh2nS+/5aRii3RJuT47qiN0Vpdxa1+Ah27D9U27Lhcx2OJxsi
yrhDIehewoEbqGCiYn1TosWb71q0t5zkR5oR5/FTK70kdghqEFg5VtprtZqQjdK1
qmURowthKquVRqFIWX47rJzV2lERT1kLdrsqdUDcMhginfI7pbxbfd24B9sVSU3D
XQ4Ktilx/dB9Qi2QyRjVzqYkpTjNXgrRwNpwixsKUbJ+6hvmLKD62m/ZYi7qWl0g
Vz1gUT4c2wDLbQf+NBB2bcmyQnBDPRvFszgiL6xwzZLUuYGiOiYRIQvF+k+ZYfrX
anpAMc1oNoDjV62SDfzLUcmHu27G6Mx4ZT9HbttO32LBZRGU/6v43wOnXqi9J1qc
uQetS66tjWnP3iUkFpd8W5m/Y0JGTdgckladm/AUyJ15V0zR4Jet3FXqppKjB6Q+
xOqKgeRA9QsuPjnxlD2IEnJw7FZ+Yzor18wnEB2AXgd7vYggKgDllhBKS8sHwnzZ
0Zjokoa8jC/LdlZybR2Y1bCehmEl3GYNQjZTSpoS4JpljaJq1p2cohxFLHYFAH54
Xmh60+j8gUjcM8QNv7rO4MEpXc4GwOLi97GUWsvqo+RsXhV3+xcg0inbUp+xanCL
Q3eplbmyb95UUuSVIchWmcTkv+w+Srm9wCozti/3W2mRkcWXmNnachFC6jcEEoDz
RZZl+wpR57Hu8WcEKrx4VUcxJhctmyfhUd2zJXUWjhYfYDu+SX/APkJYHusSB3vh
8tqflz+lDNmKA+2JitcKtE137AXT465jSzQ7qOQQTM0UdX7IwmZNrPEDObNMcA1c
K+IU5/+zfL1Ka+GeaVAAm7qQCKHq24EPLGQ1uWoAYgE3+fjzPjXRp40aycLBYy/X
RQ5zs6Qfoay/bpPPn5hX9d7x1HpXJsiBk/TouYEC3HyE4zCb+iTEyugnxWKwT9c6
vdSZzDMpoZPamIxC/ro9SZsSQF1QxjUeSayKB3J2KIkPbp3yuby0lKgVtqMi7KgQ
K6cb0T4vmC91bhZwFO/Cw1TRuyv0vIhfwFxmD+hBZN2lXw2d+EMp6HD6EO/Tl6b7
hn4s/zfNSY0QmkPJiW7gZ2ksL8oYmrkiEiHhXeyeZB3Uo4qSV1aQcu/Gn34O6pTj
BbO6Ot1Dhy74XtR1kM5Bo2yNOysad4mz2/Q/PqOGs1Ut2mR32uvzNhc+hmY4A/Cj
4Q7Pb/BgG+dYBrZnxLmAf0d6HhW3iKl+JMi+j+T2gwtNoKmm1GBWEhcZ0J6OORYh
ypL7RFdyg5UKnZrjHTQfDCqJIByJt/7GeOgDy2v7zR6OLTUPbe/h5lTwfucgjXWJ
/yruHUu48t5b2mIGvTyS5obiybPxVTseccUaf5XieHmCRcXL1i7wTGKh67NxKX13
5fd8hdKLW8sOc1hU8rrHljXMKkCrPzFLdRF+cSu/utmN+mR1EQO3LKc9km/ONuNc
KQqx/SEOuHYVoaRl0RwypNidqpV5iNKHxeFZTPIs2EbBzzbsckCh/bvUrRy65uUl
VCp7HuhiBCbqsc3TVmxry7nQ9Tg3Vk+HfkV+GCxJVZog4kvp1Wk/NsvDojEsqGqj
yIRxAc0UK6ounjUjmUew+hQiSRUbD4V0JoktD02Gr9pPbIb8nMetklrv7kxp+oQg
nX4JpcZn5jPyTz4rgFqDSKGIqH2lRm2nMXZn/pKOn1ETW9KTU80Opc5beDjjAcwv
aqe8pBfXkk/VYY3WRWZebp6j7zSV3aOGN8lZ1tBJ45pvmTB4IJD++JFevYR3c4pD
BNK7UQjOVJuBBS5rS1s8a4ZPThpGQ4pGJgOtJk+EM1Ldkeg56foOAQB765WmPrYK
x0Ez5aS60FPKMnOWO+z3xSWqzuZIGHBhZjNIuTj3z0wieKbOMU7aKRi9UbvAQEB7
H21TdQd/3+/JwFzhSoBwSu7bWUHJjGmF4B1TGeSr09uXBjgid4DqGTRVmIT7MPxz
2D45x366Q5i/h7lTe/Zu518vomxtVHU2Ny0ewSeih42uANXkh8R9N2h3krRjh5Gd
yVPeyfi9TC1ICjyB6pm0LuK33HtmQXtKlTQ4tUzsWC1g2Py/sk5K7kZMWbrFY9Si
yZ0xQlFDMw44j5hHAvplh0xAaOrJiDhdeeOFlwq6SpXPm1ovlxs98jXSALVGxdfO
MyIRD9ZGEnW5jjOR7sU2Jj8rDkvJ5hZv2dvy4ThGkZTxbjB/vcZjrkT6kPbrnCJm
a9MHiOERvqjuP3p+0Al3CduZAgNKWBUv+EIz6I+l/o6bREh6JvrS1v1Bn4/1F2oE
0QnnJ2+Ys0Msh3bADrIInGVg9xmRL+4L+tbCgsgaYLxCXx2AYbxuu8gWMs4fDljn
RgwtjQCIS9BWPtE8p3s3ezkN/ZBRXavr0g9qa7GcFVhTDnhcEhcTzzzb0HCxIZbV
gb0YE1CRWuOUUgwHR2Ce2lUMO0At8KMF1dhb9yPNuHHoIYQpVN+AchBYTooL3n4X
ISkWztUCb0Gs/f876bNO0yCbyW3ISPrF81YtwE5POzMsF2SC3GsJ5EiTkQRXFNTq
RqSOpzhllKh6AhQ8vJf8SoLmLPissTiybaWKPRPLdzenetRgRBE3UBrmnttpbfWX
WPbtV6w75HsrMWHwBZFREfKX2IApNgK2oIWp/lQEEm+mSgs0bhqcIl6NWIMTzWL3
CvEsAt0AtST/tuF0GjMFDbAltAns0IE2ThuYDxBfBwtvadbEnlAXvuOIJJg1+1Zu
uAOfcaJYdp1u1ob1+8PRui8wBL0tLmNYnOXOan+m1FbBhIggQP59XGrRwVQ/eEbX
LB//cRmtJ5igULGYnBqzAz3HMXl4tW2sEfCE+zGXVaI49RpSq7i0MdWM2jYLkycN
Mbi5G75SfBLk0Mvtr6LoYIx6acGNVVKxUPZY2RtT/ceuEyCIapvJ63iMfUDfVkYz
o/QWjejk7MS0unaZB9PY08ZN+fk4dVVDVRB6RL6E2t/PJNotjPbhZFkc+wvSetDd
hz37iKe6mXZ4stbNA6M9TjzYhVHwLTyitCPiL+5c4UWOcxX2E+ToJk/ijVnacor2
zREYzO6/Lv5zU4P0v+DN5ZTgLitSumYhO19EiZjj1ulpJYp0VE4aJ1gclb8Dnu+E
e1apd1rpaSOpMajs0cOQmsv2/XOV0OiXmzVOVmfJ/6qiaovAwVN2WHrJRYirOxSO
QB19zdvIq9diga7LOVcm3stRMg+8tWpaFOZVj6q4nNXVxg0yDU18iIEYSOgG1Dns
FNXikvFn/ojc/w4nP6dNPpIX5r1h+YJP80Ez0itolgqpzWPCsAtCF/Yp9OB19ECm
KPcA6tyVvLUuaElQlyxomhC2xlod7OCWw2pmy99YdBSEsrf2ra0222tCeTgdBQjM
h+/Xr+1aEJKoIToIInd9j2cC48P10jNvhe/5TbiMeU4pz7OB9hGU8TzZCFlCUV7s
d06BTYo/skRagg/0axPgGwkWQaqyB7v8y83kNKyOHnh+LzPKLijqjEjHeKFwEvSj
UHmUcvWzN8+QFAf2gZnDmPnDAqZMHrJAy9it0De/ml0ofwl93ARYfYks5C6eBvNa
EM340NAozGhALfGIxdJU2U9VlwVnTtggSsJa9cOHEG8MUYc7P3diUebc9DAMl6+o
98gxJFzas6I4y65oOm6C0eWfM4Z5WTtoHa3oiW29Joy9R94eKmWqGmparKkdTCpw
1chSk4ky3n3hQEID/+/59Mn/68j94QpW+PvHFm1zWlGYxkuVqr/d0hV/0s74Tfw+
e2wP2YgqxkcFtcZyRvhnAbUlh0UojkOX5xu2+gNEj9iVSjNFMLXsHwSVWCdhUNmH
PltIBnUcdE6dLJwksq7o11cFHz/jULIPXlA4WObtTGvAwtt9c2y2g7dAaAvwGoJJ
cSLKRK9QjnqHJ69o4tNpEyjWeILnoxy+GtByLG0DJMjmlhJF+yKomLx0jCHKqtr8
0j+qGRS6WzeavdNRfeoNR4ML2E5pwZzpGCCy4EYUGBMC1iTnjODd6/pj2mDKck65
pTjbrPybcBrgr/C3pjf9BTsmuQBM1DNnj9T6WdC5HdEZw4bU2urq87eBslG0a0Ux
G7M7LH1hUAwPZC27fnTgVaPtkd4Q0l3x9pbB4NXv5O5EJOu8PwOXx0zqejB1L1ok
5C9chjwR5tJOq9z+q49YwVc/INw47KIJ1137Q9SvTmFCLJXgaE1v2JkR2n6cT88Y
yR7xWNa2wWz6BXEzVY10I+7C1f1sIaEyg3kzay/xm+f6kWE+NSYfojg32o2MPLPc
5r5QfQtGMmPYL7VyDYnvN+gpuedWzy5gke6ERx5BmF0/4ns5WpGDP6edORa/2/On
18NiI41hulTGJhZu3jd3XDjCsBWXFE6LEs9QWWUIvraFJRLJLv+IALQcQs6rxyTm
Z0TK7BniOAKWiFAtvEmpK5xJyRM18MwpM46v3YfWGOk+zj5FEOfY4UnOlWNA9bYR
ughAb//wnRdDk1pU14MSR4TXqg634x9QqDn33c3raaj+CkkrBIFJQ5MIYwMTY9uk
nq2aKi6PeA1xBJnMhMIRuO2drAbJbVpmKQp6oaaR9XiWBG71YwBUaF4VzdDIm9Cq
cy4Cx4mMNd1jhMLx8ymTo6ykI/c7ZOMSMhovj1rFiKcqHV5fNaV6SFcl1FGjj//G
NimHAJxblrYXmK0kKaHIM8izkhS7LlIZ2/ZxODP9zs5/w4A5Czg29zVuWINze7u4
eRSSz2GXmAim5cVOFxtScBAg6ibqPOIB/HloL8obBhsBcgNWTFTrPk3mYr3iYak8
IY8lMm23MqNXHs7QUyQeJA0doj5k6mlRU8y+abtn0NIeVhGniM4DuWxpvTsJjefc
Vfb+l9/wfqF2JvT0nBlO2Xv+OvrSdHCowcz4pgfTfgA4/bRpTRjVKetPW5IH3FEl
xgpFb6hDqKyKYuXGsek9wP9/soQFtLM7ZKAcK9GEWg4+ti02SEmy52R8AgFK6gg2
oYA7435GuW5nJwpHwTBFegYZDIs8YmUwWxZUvYRVd9WAcd/ukFvXmwqKGxgR5LYt
4rYnRDiZAQSVE5Wl0Tm5unUlzC2ODx87Wo6a+eMyFavCWZ008kHQaO9ceUPtjwwt
RWrVWJkz5nbVjK0MFvQDyvg61ZNajEdB29oVomiuSxI7EbUJoH3jlCjqbMPofy0m
CeOgl9/gbIGxhR57vNEpj5EtbTWvr5Fy2igzSqUnFEbG0NEHx8aNNF/NkAvgrPNE
kF81YOFmhCngX8lg90iJt5ymGZFw8uD17/BJ411ZFBpo9mTvF785lcFwvbgYnAWE
jMeAPU1hM6P8eVZa+kt3tgbuSfpziXnciJDh8rK6yQXYzWwV6C8/nTLSEZUqm6nq
OYOD5NGcyEV3vnN4+Hahlbg52VZU5QiqBagqXJZtytbnw0Z7ZcWwclJqFlss6V+P
3mBFRMBGMChYTrZqmSYKDkvL5+RcH1zpHVg43o6H8b7lbtzDRLJUmXiB2Xzu0fpA
dUTb1Jy3qUQ+qsFecQbKKw7QoMlzWMhwzKTuzFUNL0TK2iJbJI+XwmMPzYfSPLkW
I5JAMoC6sCrsPIEGmpGTB0vTb9ULatBP6W5xBwLPQ5e1T5Cn54A+jDNZDdJyqCSM
4W2sChTefw4w3Vxc0xQYvb4TGE4yga+ZGC7phBxuBSBELehLpI1ka4/rRhVClkXO
cavBTAJ1DuL+xBVclMm5lghSigSdF5wS1BM9Yb+ZaYDjtnD5hyW8o7flD9MT93Yx
D3b3E3Y4kWVbjlHWr4T6kFWODHyWKebcTMBu95HLzoyKzcJeudQkjGwDrBzmVyRI
1g44Vgwf4SLYHB6Yv8ENtxa0JOjW1dvD1s92Eaxpws9wAD+izKVjIFRNv2Zhq4pL
0RpZbQyVilLiKLO8O5ZQY1UxxCUc0qAszrFqeHpmrAJ3hJ+x7+/pbUjHxIVa9w9V
AaOYi/vyp5lruRIk5+CjY3hCEnIE8ZQisWerdhZ34AGPBljT+YH/bMNtrRnQK6Ob
qfrwks1J5W7brPVzthUp5tOL6CFYFgW+M6Cq0DFZcNMmgvClPOdxLcSRLJQ9eh7u
h5ax14uuigkdI0P0ZEbGDpycGQz3y8QYNKKfmT3igGPhLe92YyiiJwI/sy0iZzDL
PpS1OpQyb3I30Y2SfD7l7zoeLNgxoZZMj3I/HPEJ3sRcmIjgVZvCjTGSulsXR8FA
M7+G/ne/xSW6LXkgIF/gR0O4WSoy4gVb/9F1JaQRjISZQqTjxXscBkNvfcTLR8fZ
Ay2MHgJU4bxqbDH9H4z8Og1/3lxtRRcyEspUC6/wM+DxsGNQ/Z0JBVVYz6hXMCG0
Y716Px1l3tYLaenBhr+MFqIbDkYmeR1QNQK+Pzteme+ZOWbB2CiF3GNPzjvYUHjl
TChnML1IoXzq/330rX67e3N+FKzyLpJoxQuL9tuxE9HeuZ/RfJx51+vVyxR8twO3
IkFAlFRdzCzMj+YT+VJ+o9djBuUYiCfClQARbNEV9ABMaCcx4Juha51xJHwKFYH4
SoU22WNw1jLLY2D1uG4DpZe4m6IFSDhyH9L7tG1q/C9+SsLZRpLP70t1tIgjuBqC
ScQBqJazB7+dlGKd6CQAXWWiCi7ox2vyzg4Nuw3x2lBpgnBHFE6aLh951N9kZoh/
w/n815gT8TsT3n9ZFnxz8eymBnL34U35WcxKhpXC+WaTM2c2JyOqeUe1iKO0C4Ez
tJrb7/2WxlGOPdk71kicUXF3qi6oh85Y1LhYWVb7LtUXCd8Wn7WXS/rgyohSRAY/
VYX/gbS9LPWSXidzQRiotX9I/l2u23kWUZTJB9cX7AaBoH4sjLXdSAUEINsL0ulD
bcQnCmm157wSLJEW3TSH6WyGWMx5jtfL7sV/jnqfhGDO2KWxtgRVS39qL/HYJWkE
zLapCOIN5V1zAMpNltq648lVYVHdjaS+haTU2cGqh2qXeL8OblSvnK60vEzKQ/5Q
mKBqcXgOvV1r2vk47WljxOlRtibcefw+kpTY9OlaF4CSvvzRm9gqzAKs/eVbQqHD
o1lfqFXyKpVV1c+zlFh4Iz48P+r3zeYjOG5p83MHqlzSbFkWranRIgD7gIQ6Fe6a
WVZ3qQ/SDuiiEgVJpFyBYNpFDD1p/02mReEAy5P0rRTDTEe4y1DBoqKXWUGh1zoX
M6n8Ylp36DZG3QtQdumkkYH15IUfz5uxARqktHaPHkYI1YEJmtKOODEdEcPg06Sa
bxoxndlRK8is4W8JuUDp02PlfOokeyO3qcz19TGgIwfhnl0LrEI6uHG2HWBicbxO
ItyZhg5vUNRvEkrW6O1qqEtaXB2qBFIBZknfJFl/Y1W6xrLmcVIt0TChDSbf0v7H
I+sq021ECR/L1ZkqZsS1md6DYRRbsz17c00dBEUGHO1aSk66RJCQXfAaDa7NAUDz
4DRO9ACrfE9d2a1Pjr/X9u9LJUsdHTRouuaTChJFjEFy6wz+gAgypId3dDEz1t+/
Q/WG5zZWRqJBt5Y/N6+YJiVp9NL3nPWX9CRQXsQ0sBYysEaTWEqizBoFd9HqUxQ9
LJC8W4ke6l6RvfCFCUISDLAHuCAH41dpKR43rkTiRXXNzshlhgqVNQcYyfYnPaa0
RD6hsE5rG36iHkyC10Qfcppyg72CicLBTX/+J7VBgO20Bt/byqNPUI6Y1o2Qh8EL
SoLYR/lT1D3t9uZ2rc+a3PwqtfCYIrTHgUaaX+QwkoSFhAZA7Dw3RUyfu8PzwUXg
hgubEol4UWnNPO48SJB7utfzP9ScbfiG9cO+T0STE6uoaMfvw8YSvIP3tp9UKEzW
kH0FD2MFWNE+MA507S8khIV8m754kfJOW5rQxKtPwED7xhAGd4R6DY0XueD9mTDj
9D/RlVogzYb96w2gQUweofOg8T2xLEzkXoyXejaTDriQ/LDKwqdQulQeS9Dj7a6v
kbSLzA2Vk8q8orzxlnDPTDCivFcwyqV8KimEt3c/k7OxeAAdKMmj04+JvQabHsBt
Zl5jPvP8oI/YPL0QXEkaevjZ4ON+chwAsdOKOEGIwIhncJ4iQIUi3b0Z2fH6UhM9
yi3cs33jIDHUD8Fqe37xNXm+qojRJvxSDvMfsOMboWq2y7IrofZyH13X6TQDCS/Z
mXNIhcXm2VZ+hMyIbLmGr0DgMCq8IYhmsmn/5Q3MiDox/E5deEULxg7/Wp8FhC3k
iXyFb0CrsEc42rmpBvcIbEZGmPXONEf5PBz5ORSOyQVfCulTQxAnVkPU0RHj37+l
uPewc4Kyvrjw3fhlGBRs/taFbiJ0B8Ww1sgGif+KGay7cGp7SGxW3bfe+q25TNat
AsdXgo+K6C4gBcOLQjMAtmG5N6jpq9oe1CXCfx7wnfWmmkeopMBa5sMzPjCNbs2f
fWgiQ/qOj99TC6HZvYQrALl7uxkcgsk+fA1nLOdfymWJVIPCv2kIXkOvoZgoRD/p
HDTXi7H7OqJl6TWknRBixbaY58JVpSyyO/Fex6JTM9PHcYdv64NJoEu2ZHBOFFX5
8sKJWvKkh67JVnGvYtEvA+maiWK5Hye/Wk0Qgr8YAswMoY9JsQ9t0XuNhRTWxdqk
14vKBHjT+8dBADvw/oSEsJW63UGScwGkCJP5B2hT2ls3DN0J+ikv07x3+Ubc+O2c
uVQDED9YnwORNOk/t0AeOsxIdWHw5yJ4JtdJxvNJJCbw/vcgEHzJy4kIrTL3Ft4C
VNo4aE0MkEnBLQn0o+gv+2p849uwh2LmGmwTlDZ6Y6MmgxIzT8IzEUHeKntI16wJ
0W3sCEn8HlaQsERAlgsQT9gfgEwFWEeQeI5CYaCkNtOzBT/eynV/l0WyoHqc0Ss9
kD+dlUFd563thZt6Z0iFff4EhUIZ7X3KATK6tj4DeoGN+NkvXnqlf5AG+Sua+lCQ
py/Q8eTGCsc7JUJApNRgZmdHtMa85mtoRV5JnuRf2WSCX173dzgkzHOEskF4Kq8Q
NF0bgKByZYCdTr91M7Ut5LPYzuTPmHCOB8KYect3WM0HmlSr5IuBGTgOIva8tVS6
UDes5/MSpzOT9qbitximZhDXnwv6Jwhok9+35xf6jyZPP++/jAItPC16UOJcByFy
fictwEvqt6pAC2KSENai+XX/HSQAkwSkPLt/7H+DG3fvfrInceVmoAGR/7m5xAKR
yQNSkFNQ2RC2bxRqrgHGEKVlLbIl6opJG0mt/ZRlgNFHrCDxBydzgeMrwkAuOPnW
v+fzDoFX5eunSaHTkF/pLKhyc+OIRE19VVezkXs2Cw7N8FJy5IbxV1skhU/mzx9B
wvxaia3KA1WYrJE8kLbkCZMiIM4Lt0SZPRAFUVWg5oXUrgzoaDC+YYJ5ob0c0OPg
R/dPR7ROQW3nrmQbD6iX1GXIojJJ+ZYOfYTAw0e4D0oak7EUYv+kPWgM9Tf4jB/2
nH2AMxTg+lPivgOKUvL2rWP874Gvg6WJFwiM+OrexRUjycwpobcvHuCSCeovfPOW
tqItc3jfcrm66k6FqWY0UI4aiNgc2p0FKYt7gHitncZaHpensPwZjrQN9sPWvh4z
CdO+j3yS1CU4ShMw/uazrK2dZZ4XA3tuw2M4SI3ZVzg4DFJVuvx+SPILh6PagVKV
eKaLF4Yke1rEtVJ7alRf39Mxv0/3L2BgpvJSXgnFrgpI5pKZCb6lb7QKg8LmSbGX
8QuwHon/YkJErZkknYcOMLQ+0QEzO5mGxad+8goPdS/6C+M/G8yPQJBbywGBM9ko
I5PAs9jBuwb9hDe0lDET5HckgMxp0vZRbYLfj/zxpmbBDUtYmcOlsr5AD9phHXe5
EnApSfFQvaJqnTEO+QO4g0yJ7H0BQKYLh7TSSpYDFLftUxpqTQd3UeG6704tENpd
RWCt7ql1l3BkG6NY11kqB646lhPSKkbbkWlxzrNkq1tPorfp/YsKfC6Y+zuyR7jw
Tq514WhCtGNrd6ABn8NoQB7pY9wblVGFfnAk6LIH2sUOnPQmYZ1uxki+siV/vFbK
JrTFmk4Wutu4bInTCJl/dRswvFIPE9C4cdWBiEaxMh+Ia466dIUg03bYJDN9X6lw
VjXE6Rs8LPZOdOS/ic2loBxtZWonH/4cj1fzize2GIauWjr+ZtGuWMvN8f57dwS0
MAFDUhKKOiWSlU1YiLw6f/x7vXLfEKBY4sWsDBOGjPLQ06rsmOe7e90LdMoh0eQG
fNUeSXB/JMYjHfy5knM1ntp0PVlfuNcdeTCrawiI1iI2jmlAnjSJBJ9n+PCc8t4y
5zsFf0eQIqjesUhZoJoWlaSUafTWxZS9LerPcqzzzx3PmzwWPmGfG0YUwWUv8P0D
Xto3G2CVzXeYf9dvCleq9guAn0TKSJQJLsWO9IJoAWs5XaY5VEWJwcruyBYcSuG3
U06pqSk7lifeUAl4c+wQMu5vPa79Rypr7rP8vwJ+29TOQ9S3p3O3jT8wGTIwstD+
gCeNs13t/6MS2+K8UjBHNnsGAfIBAuezSiY2nRpGXajmQzVkUTt4aZkX1ijn0ibb
m6rug5pbwFy/MWagQEdxdl+DSDeL/uSIwXVto0hxj+80/nbdG858HQJI3sye9j9M
EWotin3nbGRXKGVWjLDdMn/YupaG1cfLL+dYI746WogGv0qJpjkd8f3m9gDWqM/A
lHVeERFYfywTerZ61rd+3BsIzZQtyuaM7MLZrH0MQ6sgjWJjjtlX0xMpF3JWwVk/
tZyPIr+jBrFCPwJgYDLRFqiUNyQMSFXuJySxUTG7DjlEiI7L16TUvcz1VqeaD/se
8yVAbaJXJ1gecRLhXWuoNstnZafa8XZJ0mwrlsXHdpULj1YaSl0QKxuVIll+4foL
JHoRYzr9iRC9q5sRv8rHth27SWVcUjRGep+W+Ni2T3T5SouxddeIf6UntkaMGXRX
Ai+6XALmIbZmCACOaPIkYFURSl6JX6vX39CPtQrMsjwfsdmiWufaMcLLlUGNVA89
ahr5JBM6dQ2nV+uwZ6ul1eEsS1gWZBCgQYGWLXDAeDJLPlFId5BoPRcfAs9QiExs
Z2Q78O1rzvG1uc8bOkfA5wFnkzfLQuAmFtJ6T/H4GvPNJ/Sfvvp1NFIuYvkNttia
FLuznZnEQHSMdRz2rJL6M/2SxcuykjniDvC4HXqj6fKdbSJsff24ELEJpwYtkJQ5
yoAiIO5wq25l8KqCcrqrRkBUyngCDSJBD/n37vpqnQcUqzJMCSoIcxfKjbikrhaV
58QbgLZkNYBN98pzC8qF6qLVoLu/AE+BkwvuG8aHMPC/i/vA7+Lqzh+QDH1czz7Q
RvBPJ4EiOw+xJgpPYnM/CLMdu4ymDgXC7SsZ0ZvH9osIplaanah+sI1Q3OjI+4E5
cGqsa1oItvqrQeNfsbgkGwcaMWtxxgrmrJwbwfnRHkIfRR8VbfctfLi/smZVZzpY
a3BCBQhqpnKqgPW7QXgJzmxkWVK/hx8Zr+xcOogOiOfIOd4SyWpbKLNfsmeXZaXs
5Tir2x8ILv8rQkxU63jTxKYgeN8Nu4yWPMXeNYviQfTzqavEbER9Kon/EcMoYFgg
K7HtSB+rcJsQEFoQ+Xy2mIw1loRprMFu82jQr5T2RohzF8j9CUbz33xKIn3mfUc6
w3+z5+RvNOFNNS2GGsmsYY1NPM7hivnK2kEsNPHymMPmePz8Z3w4BDBcIzxF96T+
VOcgRbJpOEfSFYfZvWddIz080wP2d3d159I9q+FXICcuk0Z8jDnZQcFG6dEvA3J1
mZK5F4ANxB9Ucs/n5sFDeDNrEV8epiwmErgprvKdBw/8kVo//d2vwrFWL0RPu11k
TFb0YpkuVzY7Q2NXO8KU3665jcoTX0axsJYoqp6QWPxP1CnNgxYnu75cRpNB08Bb
jZX+cPj5Z5GFwtYqyTI+ooVx/h36IiYkJzPIKV4AhKWJjoDiGx9RrTv3IV99TjBg
bgSxsQ0AYApkHINHwt01nzyLQszVSn9qqPOzzz4aiBCci4YljJQSvBQJzcH0dwUP
u4bZIJ5zYtAqf+4cv7BwjH3yfZxy3zPGxk5+8NOsFsy6OVcehJXd6T8xGgnYkVGS
calCjPhTn3WtBnC1JNmK1Dwo8seaw0fFGAWxNTmJ1wWXvUzPJu+cAAisJP7mNwOg
eH/402InBJKwAX6XV4wUgf/3ifbzXVZSY2eC6mwxprGkH6Z8YwZjluJF6tMTsUVQ
ET7KnvsnpAFxE6sGCiPWsKE/n0+DCDwONQF9N+L1J5j4kL8XQyLZMq1W9mCjY9ap
XdKKGzav7gHG3M9FYNKo/+FK2ludpSqEUelYzSvrrwse+Nwe71gq6aaQHUa+l47C
/c51Fnj+RyJ5Fvi6cvNMrjRBNIdblr4UhnHZBwWW8OaScINKm5lBFiTGdeptBmjm
8xmTkyB4ME1nsS/5hUE27K/petNztOf+IF/Ga+JHgmnl6kibVhKEtQJYpkuLzu0b
waRTvkT/obx0UJ/uHBHJOjUi4N+vKCs7xTui88duY/Th96nrEL5Tf39eo3oNsk9C
/Q2xDf/Pv/RapSzpATZSOcqkvysWU2NP9rAlkG6RxDPr+CgwXUG+G/h64o4O02mL
bfCppuotK7ysSVEBgSJowqSPhQ4CaacdnIv2jcVToV58+kW1N44CVPXlP3Yax9Z+
yU8UgezWqL8EWToFGkyYZP/HUFlFM7EaSTrAGbM5Rbdh5cZ+BXuSlTMCihApVHnQ
60e3/EYaVc0drUi7mGDmEWiz9kx1XBqJLBLWTLEk7CPoNICI1Vjejh5tJEj+OPVp
971oHxf4QTSc1HVqtdP2RL7nv5bEi6HIyThQvv/nvNmqwaBw+feR9fFCizJxvPtw
5lRZhecD4rSLOV+83+LCoTtaZQhGUQHjA4zL/5gVUc7mI9QO2Z0kOavESVaVYsED
HNMlJfTg/Kvo9mOspfioIlwunPcSroRa2+m+DVk27wsigrNZGPqQ4Y3ASB7PrhtR
03MB6WPuDxA5Y2tYcQZo6PtXTMNOUYa4jlhY/+4wriwA4USWNh8Vps8Zr214WTu7
X7N4YggSaHFQ7tih7ytBkbEzJ9jdvX8lr3XE3McL2hqq2I10uaGP1HmrsEL2OUkW
CmkNSvqQxvlkBEhsZIlywKXDQIYLCbHX5G6QjtQ7sGVemU0mEH2RF1EtCxhASOeg
rpjX+xlmJHMoRExYdHFlIVlVmbWGLJU4JrebVevABgnLIwlyN6pp1c0qCMhXL5gn
clIpd7rE9v80OloENSGcwIFmZOFDoJQMasjBHMh8gMScfcEt4xgNukOekJIFIYZh
BGS22zdLgeb7HfYp2NbRpBo5NRzKj259XcyEaXNM6iBMkpMVVy8Yx6zQ7JPWTLKC
ViSII1cojDXG8gX/AZDXQoi3FewLNbCfNuiwPgK/uVHRElny6EVAkTSTB+besEHJ
pCxb8x/YcBW3Y8VSHfLkGwzdp/jvIMBEA9lw6M/C608uBDuMULIhznbsvpOX/38b
IDNDHs5j9rhNNt9G2VyQfVJ5YCXqVMtzFeWbfpQ1UWhSR4NDfA8qhn6beQb9fAUo
pstyQY8AYXW3AFE9/6BxqnNNkxesAFRx4UkSdXNyM8IwAu48Jwzo3ItO3elLj35C
/BoCyJeBEEgU49h3c74NcjaYDOc9njpo4ujTOwLcNtTKsCMEJ+jxM0dkEeVpNbIE
9KDfOsGVQoOMjJ53iNFuZDbHXlpw3A482h5CYVvni/IiDOCTqAvucKJKwswlX6MT
Qb0kVvRXr8XKFmrG9iV0nVh1DraprHnrTUCAYLjmQ6wfD1JFfPjzW5j+0eRRuvj/
pULNLnHmHa9DoWmTF0X9NVyqHr1Xc8bf4YUA0Fe2YUyPGZjN5nW2oMdmB2E0P7MX
6BS3vMq/ytGMIJJK+MEFnQGurMspeZNIn2E6u/E+4cxp/UKGyD2GecW8pafjtmr3
Gmaq0s4G+G2bS+4pDrt93G2OvSJFqI1PRfhdyN9zJZ2Tt04mVqFEJbeB12uUGOuy
Ah7dIotBRFSCuhoKO9Zu2nB/kk2H3ygZq+aGd2NCdNIEqW1Lo/0MeVmpHuO2AnBo
WYuNJsVJ7XRZeBkYHYGo1tUueziCzMg5L8z8YgWf9XsRmRHYk+YT+AwbmWaBK5md
bMRThkdXB5ly5onzgJjWObMOfziSzcbnVnSj0T/+SCvYat5AAktoupMfFP0NTSnz
h9UlpSeFx0mOSJIi6uhnSsSPEHdFhXKaTBQmXF4Tbeyp1oGsI2yjTJRSxY0yToIu
rKbmRuDTafXR+zpS7vT6R6Qhrur1Nt29Dx+x+wZw/VYkfdPdcQP+3oH+GC9TIHx9
3DIXkbXIZiSCiyvB9MadTBTFl4E4HGFJcAQaMpxiH9+kk/9aY2tXFwi6vPEalUjj
FqrcLej8/hqa4hM4srKpyrDE7p4KB3od7mM1tFl8GTrNZtt5NBlrBnABqtW1QeDU
g+MuQ/UtbOoayQYmptXdae5KcGVE8luUadlqLpWUGORS7e5DICLtt6nCFPT2Sw7k
awAD6fi539kpvn0MBv/cZr3/DY/FIzmC2IIbLr/BZKiPHT8bI5SzAcS1lSh/pr8z
WeawtdHJ1HB1eLcGMpC9vaKrFEltz+WJci5wqzHqfLvM4JHe0r80uEtqNSrmx7lo
t2Htlj/z3VEYnjc4gte3y0wukLuvkw5LLxJtGQY0VJNHVtUtMuxcXNZyhknx9Im/
jkb3aCgp74aSP2x9Yc8BXA0jNyxIM+4EQwbwAChgL/pAHcpl5XVffwH33knJH/L7
GOf313ckygQh5lzxyydEnMqQDvTTe7Md+wwxpK3kBvW53GPOLVnhytZFxeTuGOqp
zBLsXPhd+FNuShxPDFOQ/5DJ1mAlLReWNXq9G8p79FWPff4ylXfNzgulYzMFrRsb
ZK2wIOuej5x4v7TYQ33B6CjV5k2Jl1+TqsCGcwarWJAFYeDPpjucco0k4vNFbHpR
gdNt/0KlzDMik+ykSKedGKmOZsO0PjZNuytRoSnOd5F0fU06VTrAmc0OXWvZjNlL
cf9nij1Gk0S/T2v7c74xsuYweAx8Ib7z5N1nh+8Z1i6Ii4ql6tmX0P0zlGsHPii7
3kiAgBo5jflv8uPTE5bxgKqcH9UIhwcPIhpOtIDwUZXddByYaO6ysv5Obx4TYnEv
RoDiIOuNPW+dIlYjtLvGgUQSyvTbq50ril5I+SnDRuRF1zZvpuEBhcldQQPOIYce
f6UuGVwSs0+t9iduCozo2N5AWB948SVEmTpPBBtHbjctpmnlvR2uO3j7OVZwKlbZ
mV/LmY/TuzpXdIIUn2tLufx3bVJoe/bQwnZDb6HGCJE2FYqeyVu+dzJ3vTzgKGcD
KHTxZV1by4jqC/YMcO0A9pOwfO3/7TCxSviIZDKUL1goKZtAtAsjddN68EN9grdw
yNFqLZOUDD7NkpNN59WJCbx7IX6ML5CvBE5NxvWL+/wmP7C+3nUrNZ6GihLvSDiT
XzOWatgum5S0xEF3k48PVpe78y1JWvXS/qgOWBUK2TcZ4pKhUIoPbpbLieyTyOis
l4jRQda8s1+i1M7ULqNjkIJc+rgEYxM4WcTu5ApkQnzWTVZz9PcqrNK02y73NXnx
wCTzkfeKVeoK331InXctakycVlEh5NlMW4VYu4JkcbTs4gDxMnY5d7XZJV30k8F8
N4TaKXCIkwjr9kHFZsfFjCphyjhyXg1UyrsZWmR8ThfcE+4hXuj1JGwn0Qsfo3uN
RvbpQ+bKDSFrZYDVlYCTUHtp90SNIKcoVJ2rJCMHtLz+iSdl5AoHP6TlpG/tnc+Q
v5G9O7I7i42B3d635GS5v50/b4rMexFVDwKh/V0gJTMb/yIAPu1HPbc2nlcyPulu
HbdHtt0rZkSuZKdQyi67fCAW0GAJiOqTRn9OVR5MCmAzPEVuVSgd/sbG4QhmQ8FZ
/ckpeFFWGn4N6hGiiTtTPNFf+c8PcM0ShwBK66x0FrOE8s2EcLbpErUJa7r1yuHW
zr8ywneJ8F5guSuVw6ttQYWS3QJnQMQLWCkdy/31n8mIZp8zj+tS7qmdurJyE/VM
eeWvjt58j6kAbbQqv4XB3iydN/TVOguPsuO9/yeYJvNhHFDPAd59rJ8nMlgUZcyX
925l+nhrW21b1zL9okRjjqow/CErewf0AtGpQUAaSkM7f/zjEneeaXVau1P1wuRI
ppPh539th+vhFRaJMhfWzmHJHpEDotvHRR6uDB+rTgZXfw7blM/61N7bMCeLZnHU
fD2EtpampnScxOSCPq5hjAWNGdn0o/YZv1cjoMKZiK7DRSeuuyKnFhYR3Q+y5dIj
1IuPD/bUl6AiDWSrS1nnEcSZBMWiCOwGRvUpNvJPyFc39brHEIE4VZTvrYJrmrEB
RiNL1vuUvdvd9yT2HvIo3iwV7w3Xn16A2kbsefBeJgue6UDnnmUIEp8M4MLqMxna
nuWp7G2h033sOVB6AUvfEc8dpdZCts8E8K3GrZN4P7IYkMtwVKvv89Jv+vwxtuyU
SUCyVVvlQSNfsPBTR2ThqIy+8EVoDKlEk5p/+wCzmsiAwI1mUr2i0ULP5oaQc2GN
HchgcdhUl5oYGo2r/7SMNxe3AkajyohW+LrPKorHgcQGuNkYYoQKYRRoFNXj1KDh
4KSTrdRZKLPpbCmItoO/UlB/RYTr+a2OUSauEJdVXUFDfz6SWNTDt+dKi6pWExHQ
1QGIlVAADLFy+MRpVSqpTKivj89jQe5I9wrNUffLEPjSBz8kPBem8mmCSaIfGlex
y1iaaOQnyYuYJW3nAivSU72c2X8xhWBR2RxQ7NgHWFNI1KcAqNw3OZSakddipJFA
2LSNjtqbKDQDwLoY/NPia+bnzSYisSoK2w+pCal/XzFsu61hUSrgTr2C2xEfwSqB
2XEcQVQ3pUDQE2WFJirxAJzrVLpKor6W/qZPRLVjnGFI4+aIreJRyD+mUSwb9Ft6
/ql0gvwJMAec7ucpRlxFEqTwbiofuRCZLJvIflbVHOc+2ir50eA+jXZchGY+2gQl
V/hqWymlJHWwuWV4/n5u0uC7U8fSt967ioN4ovT9r+QKEQzn6V/SeCkljFs6433K
dJF2i2sn65iXhII0uYJvCQN8DL2bHl2s9/wYV3BIgMfc2asMde5YQe/EjLlqujJV
GCWZgIWEs9f6M/mUggz5J0rOxV8TkHQkpV+1rv9MyrUNqm35SGWVxPM6ruI7y0a+
OOmU+UfCK5zHlXFukE3cUVrhdZ74ucO8HZHaCwP0RHAAN0HoL75HipcQjLvCuweX
lu7Vp7Adwuty8J8Iv2LMfFUzzJHIuGMGoH8WXVA36JxSQbcw6hygahi/OBr09/51
hqfqYwXw2HdhvzPvxOKtUYca1SnkSQ/cbYxPA49vpzugoT1egk45rdaZqOMY6yAG
xFNOLoj2wmmtSTEd5VAlcryWEM8TwV+mSOec6vVHxltk+Dt+NveXP3uI9GemS3ko
3gPs33WRWmODA1+sXvdM0fcBWkEltI6atGkbUUudsaqIpwuNLBLiwnXXSMgbnulW
4DgEZIq2u5RlvS9iYLVrzG9T6Bg9UlXstimiys9RkEDSKK2TpBKidz+ebOPOr2YI
V3dptjkjva/zEx//Ei7R0XvZV/QoeK0ZUos1wYJpMnfD30wdHiUpeMLxWqMq1qBj
jbKZdB2++zQZMtYHoc0FhE04k/jW2dwUbEX/ZiBtMEaGuoXpNOrKqY9AmFGj2JqB
HbpXuaaNkmVMaiFJEGSINEgKh+Smi6FAJTlF2bEzOIEpq+JwYmMN2D3eA/xOYI2s
g5K1u6ruW0K0kT7B+NjbmlpRxqwEY9H8CBYEZhdBdaBTAq5nz1V3aUzEZYo8auVd
6LCII3y8QSBxA1KYeTc+670F+lWrq/1ZYRaauOKce5fmMf8rQgsq4rXGnyNOS3Lw
C97RYXm6OKSO7SNGqV/IeQqPU+/fmGBI8CEC14DhiquPxH20b4ztHO86QzlhWr2P
/zBFKDzOG291H2QlqP/5LdwrF6ZHVIiYb5q6IMkwhvbHBUFzleQTg6yKPuVr15L/
PO+G42uIaDqqbK6ojmLL2DlAJD1DRoZOUl9pOotDmlu+JJzxPQvfY6eAu3HEv2FU
wccjtblJsTU0ioTBW+LRZ8Bzxj4AXOsRmRt84e83V4hWIjuNBECD9A/bR2lINmst
uN0BCayHyli/4mdAdGu/AFNAZswmGjZUHtPLi6eoQBl3Wl5egoP1RrRJizh+3meX
RR+opS6EqrUJirISIG+O8rKY+lvfqa9QEdpn8XdzwBLBz68YcwfoBi1uMPXI8U+f
5BTW/q5SRLrb8kXLYMjTSJ26t743mirFNJPzKylYJNCKlCrivTSwDhQiTVJqy38P
zx9iWRRTfbnw4zkBifuZ05A2BLy9BSpcZ5dU4mN22cd2ajjzt7DhcGk8uTPh6Fii
aVYjjsxUjEcy2C+ZBCdWGKlbqryLj5DlrfNODh5c76XOKXFUo9lFviYKVfPix3Qz
scowlAW8L+QmQumtlsjzKDwG1uo7eyKB3/P+qdOahlSqT0zLgn6LIJnxwFFlm41R
Hj/b12M6GRIY0c9MtFTHS2CD0tTnSb+egGR7pH6x6VmCIROSCcjQUC+SQ22ebCkz
oGHb1k9isV3YKtvjRu3SsdyvR0DGjuLMYZku7d5/IUV5mneXhAIk97+AfkIFpGJ3
vXsvGqIN+4JxQvUoz8kvOMtGXwUDNrdtLnhl8LxJcIwqspeTZ17PEyQ9yQ2W9A1y
PDa4reaxoUlJtRpovMpg4VG+lk3G/i+Qol6E0s4UHnQ+fTd1azfPAGu4hepkL+vh
D1Nc0Nx8pGRO8vV7oRysvEOQLemFyEGXK4/UYeqSQRGN9cNlgjS6e0Fixr8kjC8g
OtaA8Yh+vJh1Defqxi3GXHKCZBqPkpV+iEGk1cNGm4mDnvEU7xykkyeA1AlRkSI2
U/1uU32A05k0iu2pLD1PB3UewF2n60s8zbpq9vU6GLgOlKZ/7Ij8b/onRDjwZW33
/Y8fpGUcxptlzc6xATA7VBIPkVcPoTRKb8dOzy5t7OBwK3XmeNrqcRwwzZq2ggnh
FXFBn/LSGYkA0wPib0ze+0N2RAfcH36Zx0ZyT81LRKAt6Zlh28+qEBHs7UZuE2vH
euus8uwoGFvUuAMAlvNLr674ujK4n29eFTbLL1yvgbJQd+8TI2gbk68D1ahhjupr
hnMtXZ6Ozwi6OjriqxPcDRH2xCrJl4rDZCg9DsBe3JgvAHcdP6FEyCSKMCHIYl23
hEnW4fFQ3Y+U3YZYEMHea4qdmFAiJnY/E94MC8larAWTbDPgRURwyXfayNiJhc6E
SXDRIvAX9yUMsgDjs2QsY5w4qxiYdZakLSpbALcaN2eeW1Cf4lLLsIXn/JQ92lWp
b7+v4Yj7znoE7gTtLhpaH4IVK/zLLNw6jQ4++g5W7AxDQ4yogmjmkKwvZFnrx/gE
C/dxELQ+RTaMvAhtZcBLZDFLynBjIJxFDRXy8CAvcrunX57e+mw9JK0hVHGvHQLE
VJJ3Jcc8a4ubfAe6FtuRFM01dfryyaqYySwVnkvmngDpRFEC++H5W6aOqpqmw2au
vpt/2ISNq8gz1gS6MzAecT57QERhTpweGsaXKThQxom5i/3qMhapZ0F726SiVzWn
8ifTukOt778THYqMYv7HeFMUznPxdH8GDlCQrbOkbTGuWu3c6pRuwosdWry8I9Qr
EvX66vEAIZQegUP9aXlHhHpyxnuLCjH6NAgzoH4PE/8tl1A1+fVINxUcubvh7sWb
/e/XQH3HOmlnUmiVNYCt7XyWSgHq78qabRit4g7CKGZsCTNv3TP05/9RT8oKhANh
sTARK7oz7UhRc1JZcHE1lMqCNtNZGSj+Vc9Wl3NtHtMbBp6i6f2CLCNKFWy4Zdws
2U2Zp2DIt+UZ8qCRjzAOQopYa/X5Snu7hdPG8UJOpYh0k8Bg0dEZfX8Z4RmMBdaE
p01f3nmfVdkjIuTiudXMIXPFpNTLnZUBjAWHdb8uIljO4L5qGM8pmp3ZDTsOsKVh
W4TXN9JqV/M+jK3tIjS3v4JZQO8EgM9c4t1u4rtC5Lafbn1udmWNQa3IFlyAhY+1
wGsWmBKKw6bhoAXdmTuGiJKVrA0FglPOW07Sg31M3m92J1X4nA/URbLfhrlRo5QX
JotvNsG1Z0y4bp8etuT7qESnVnWnDDR/nk8tIbraQfA+oZMYPRxd1kPxDRSgCctJ
JsFODaBZJimkmZv2qqIGnMrhrIPOakRQkXEKu587gfCsPSZPejrtCXY5dglAjfCh
Z/fZNZl1rnb/iruIVihpmWfhQRprtqE/psou3UWyZugJX16OGewBxpgJMr16jQ2a
/ZggGM6tWf+4UJ05OibmExyMT6XmTmA7Hw9JgKA0seW0FUP+ubAWUuEojdpG8a59
QCqPVcgix4o/22iGONpMeKkjtH8u3aOJ8T81sKdC1JgzNi9i1rWdgsfSEAOjzMgw
kiHQjpRV1KTelRicIuAV9xN3uOC7WBpb4dHk6aTOoYv5rY23EicRS8pKzJ22H377
eOgknmgNbtsO0OHMLw2GMYn5IkJCkgLRg6T4TbvmTjzlGAh3hmG9Ld+Jok8glg6J
umKqEJfcCnMo0LSTUHYqnHSbkTOmBVjpHeRqQ3AdP/KiA4xwbkFE6+IOdz7hgmae
mS4Pu2i9dS8Cr+uZH1HoQPXMq526zXjG3jA/1jxqHMl8yaU1ms3eR2MKg+IbI6Tx
dBlaABjhz7D2CFHNxV+NuV5ifWaFINPyN2kkJjfvqXOJ5ykaqO6fDA8RVHVm7i/D
9mHGmHx0p1w10Imccp220vAaQmYcRPebwz9Vs+g81Cao7Yk3CXuwoLCG9FIWnT9e
T54Zy6R58YlCwJv8ykwMA0h0ptUpnPMZwM6TV1tI1KhfXWNeW0hB2fYt+aa7jBMm
Ah1wa4mZwnrhhIfz52m4qbqHV+ZpDvy9Vz5cjMdHdHu+3RYZURx64aQksRbEdjbQ
mDB6ntB+4Tyox8RhfFNMt2EkjJ6hOZYZv6V210MPjJEfxaLcC7wW2UJ9gB/cUyxb
vgLjQ+dHgCGoOq6ligDLsTT+auutgn1bW6WcEqDxdrgHockfbc55yeC44eypuzMZ
iVAjt5nEE8QLhvLvJNgWdOMqIr/dDgTFLY+gd/YZvBco9mdZALsdKP0LxvQR3qKx
U3nQIuVuf1w5u7dbI1CG2WlRg11+Xz2qyt2A0d5HjoLqunPJPUrdlQqcbTTY00e+
V+ERfBe/zClDfoB+1fywZDFDYNbPH9/V/r979pDu1KtzpT4k3asaEqJnS7K7WxKq
fDo3afZR170hnSbOr10ufGOqTOSL5YzqfWmj7H997tn2wF3TsnImlspQMyEBlqnp
sNYxalWa9SwSeyNNp3sk2SgP25/pnSvoga4mq9zEK5MGW3rOZExjIbVGGAYZg/LR
akAfKcvH6QjAZDfadHj1M/gcFT7KdzOHJqkkvoKgOoNJnqkSsyfNTf95Ak2QXxsD
HquxIUVbLgqmsNzDUe/2cxdznP8M5igdNdoakbh0yctEuLyY8g5A/8qYsAghN8BW
vDsjyGDO/315cTfTDqlzS85LGHCPp2J6/4IwU14UvM3Gtg3kUf5z0Ff1oU4ZC4Ma
1fDq/OyjAnz/M8P+pqasx40iOBjOMo0dYz1koC7QISNLZILltx8Y2Xx7f2CL+TXR
MzxhHl5SrSLA+GBhu0r/ASo7pH9f9gXNKL7b//Hlku/pxKB1z1nwuXuGA54Vk3FN
tyytXOyaUf0H0jK3+GuuX9GAvbNLxJRKRs+CoiSS9RO7j0J0MILIDfh4/ZE79p87
+EJUdEj562PsrHXaNCLcyaHm3jmOe6V1ieb7nSFfa+CS5beeSx+7P8be/xrYhB7I
WJNmtjE5zCHQ0+7vmhNmp2U4Vma5B5dGtVXVBbzWEvCqu6kroxN7oE1j+OOopqXJ
9Shcbcp5idV403nrvIsn279Mwxq5j1xNEiDgWXQobpiAq0ykvYBo+MkxzZTe1FDK
8hnYf/kyO4zEy6FPvtLmXiJTgEtTVrQVj9LOdusRAlK8YFMcx6DkKK79eVBO/wNn
xNBGUW4cJ6nSfhP2TPD7OlUlW1XdUDASfIgpLQ00lAM1RWkvXrSFBEMPPdaqqWOD
i5mxuEU1OE186Kc0sElM9SxrIR7PiMVVWkf25evJhZ//FUmvL//e12kIKh6APR0A
rUmdx3n+25mjNRjuyYAjBc2pLW7RFlkar4Q90v4IV6C4Rfs0k1RTfEtrClXMvSy6
xJ4fX7giYqNUEDc40IIOr3KMoEefDqHoEUdFxAqk3R5PEUSrU9jlwKSR8NTVh2AG
HmMfTLCcWQbzB6XLvRFvUs59FloKFAgAiZvdjM7SkU0nqewzDCnaw4JuCT7uEhU3
UHlgRxr2YrZkhTy2C2OoYvFi2o7wRVsbGVjCWQBLBMxfkHQw8fIT9UerDEAO1xY/
ulrQUR97eXaMZcX+Pr9Kyw3rp7kbJRF+hTEYN0s7FXy1ddk/zRnh05mY7Lx1o3HR
LdBecIrEGxhE052ZxN5ztNTpMax7fgTqOZJty8t5iQ+BN29TJqbO8dd1w2X5bOTU
7Fc67+EiQQZ9TEmxDZ4mHZK/WlQTbqv/ONY9HohXoj46DJ8k7ckk6X0T2eyJlrg5
P7aC1D/GaGBUqCgOeBuOFLe6A8pFVoNQzjTE6CvCGdNFoK6JogqLr46xacglLdg4
/HjdFIyPtrWOtyXJQj6lG/BL1IwnS7fO4slhPxgxAryVdyMfJ5qRyGfa904U1VDH
UcPIAaG93QVCyM5yA/YorVoSyMDyKJzZmMuHTreBmsL97lb8iaJViHmwv9ECBSlP
oeJQBekeVeGemhrAVAHtENQkPBA+rOIXZlPz2PshCptIZ+h2x/X2yjoD8NQW683q
EWiWZyIwSWvN0snRTT5OvzddW4F/1XK8kN5gt86PiM+HsXi6MtwUh/fJsVwFtxnS
Vo5jm1MfXbWL4fcctoa2vzGwryZYuTE098w5YSnmCbAk6CdIkKKdRnnVT7lp8SaK
`pragma protect end_protected
