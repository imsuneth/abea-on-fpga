// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:50 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JlmoKpAVY8iqhCDBMtI871t5WBzk3/Z69ADEeu8U0e2qjf/1EZK8oWQ/881SXFHM
9zpcs4uRRD/291ZENxGvguvtd9PQJDpPWcWNDSo7yM0/V1uXmyNjLcL7tt9lqVtw
yhU24ITnUGuLkHV3uPynDTM769MD/CqDkgnXirBJNDc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23808)
YiOZJY65Yw3MCRRNzhJXVLV5N41i2aoqjhIfc05ybHjGNMXVH40gJsolAJ7UZmSY
PluMxa00Vf/e90hel04asiaFByUee4hL0NWXHae1RNV29T3T4VUFABNsDAnaREoU
hnfZBgj6X9z3P+oFNXEpvmG/k5vP0vYofTnAs0oR4n5D3Fy5rTzz5f9T/Z2Jccce
ip1NXQxCt+ukL8Ve2Rb2VVzE5JP9x8NlCn87X8cY0ZpX6P9n+Hm25WVME6nWlFwg
YN19Wb+xheLo2DUSJEp4Kegjg8anPz2bJoPJZNgsqKWcxq4lM6Co2fKPYw/ZGokr
P/tp/1lIGaZD2487Ek+DIwq2n2DmGXs0w4eQ8QSggw/8qGeWJiPfZ1RWFkIrHUAI
Ors3vEocPfRn1i4U0M6jkeHM1HHUCBzXQmuMF8DCe7BZfegcry3CvESHG52xXFGI
dtgI0eiBKfUElLyKly02oa+18PQirxzWSIqLjKWzdPkV1G0qSMKb8NvYKdtvwnq/
gpxsjch+lAJ7OM4k0J2MI/LM5Zi+MDuGBCtWNj//S6yCJFjlMfrFRCpf9SM3uklM
YCjwKw4NJ0UMWO6qu0CNXkIqS/2O4bxcOlyCA5VL9MX3kuqs2Xx7sK8ISt7mf0oJ
TsDhXYaVWB40L6myWD7MQkfsSDBxNLk2qA3v1xl1BeI97YpzMtIu0x8agcOXmPrW
fCZtFAtKEAobVbI1L+rdj2QKI8MHhJMtW8HaecbPT9zIVDa+SBgVajW42PYgR+jw
HAUEj9y21U9JQNyoBd8lqv6l19yie5QIHsc6eOqgW8F2wsVYDtPZwdhUrDdEuXZ1
tpBkgxWFXYU3dkr1G7YzoX+qao/gvxXfOBlPuPNJtHLCbmhIcGLWepUSMTD2GPCI
qOKMpRvYB0YThePWYwfN/Cc0pfAWWR+RwuaU2v315WzQnr/K0OA4TVlex8+Jd24O
NKuz0Ajdua0VaBtxJlnvGHFsqE2e8ydEmFGjKo//FrhUoP1uEIqkSh8rO9aOKPnF
JcetrMZzF4aELh2VpNVvUjD0tv6iGorKoa+JDwu//fEN+8YOod9gYMFyWCQu0YyM
ClVmVHRnvDymlhAmXBRi23JWOyZ4j9Ue7XCYHC+9r5xilQYuiQuHHkPOMf26JN+W
qR09MuVhCKBiEnkfj6Z+DB0e6peALgfKbJYPUk89hBUztA6Y5NWOMAHwHdWGqo/B
8uk2cU8RLXCVT9c4IF1ehPQc/A/bq/tiIONc+sdN/V1fiG1bzpf3XnmdJDa8ZICB
1A3kLqoZK1ISWY12pSlFDPctxM8V50FlMBA8iFKk4MpamIoAcMkjDVkW6yJY4ewd
zPforGi5Ix9Jihb2N7uMP0J0wLARrN1hYjHh9FAgb4upLc255R725K9yAWWVAiNR
GB0iGWJz1c1CrLcZxyyH/FAT/M9Tjf8px3BCxuwYZPK9Q51sUwKUJNPqi921Q423
ubanGK+tWE1QUuMBAw0dPlUVq1UF6Q+RxiMe7nY8r9YGxPumkRyX8j6Uv4HA/RR5
+YS40b0q4VzyLZOuc8nv8KEnbKYArdOHGpdBv8bj+P3PfmNItuTy0ukh57xxnew5
vqTWKrx/T+9lORGrFj2B74Y2f55hp1d01q4aLMUgy7iNoq/22ezFMe2iUrcov6Ni
t4jMLOrCfWSVB9x4YTF3yfujb7gCuZocdiCV8a2UrIvFwJmlRUTZGAykuMXFyCcn
zr5mBLndghWA4jJQekfgPbJ1wZdHhUAQYvjBPXkve3p8FI6bCL1HNmjFNzXLsD79
+q0tlJtClFn0u7Ln1YveMA0S6rDhBaR18MUZd0fcCTbOxYfsZhIi4CGd6HmfTCPv
LZ537ia+diMmvSFkcf/2zUrhpcZlDx7yG+sks++BQG3mbK2K2gPW5107PY3M1YOp
jf2GZfWYJQ9SJ0WsG7okJ9oaJ/qdAGIXHARZ0CdU5w78qj93gxJssoeE2syyKkMa
xH3ngjvSKJNvjU5y5+eJPnt2AoMLY46SL69mLSYBXvPIuttNpDOCGcQqzA5tuEfM
Nk833R3864cDW295kQP00WD3ZwqFpEERDOGxJ+S86Hfiai1tLyoahRxrgpf75RZt
Z5dWMFyvWPbLuq40SWokEUusS9opO1K6UQmyHsNrIv8OHgFFXLLIAEKJpxjPgW+d
mtihCzcBQphl4YANhJUVMvYK1lgb7uGzHn4Up5vt56HRXyc7l7vPA3LQUWkmAwzp
WBP1cdDGBctNMuQl0ummp0L2ozOZoW8PCveTGLrvg8LIspsbOHMw1BSsOmhXVvFd
hqQlnAGavFIWmcojrK0HdmJtif+5JNtLkrzYZmGYfNLbTmnpQMFQ5/cF/wscEr+O
9CQ96HX+BHjVmUsY7ipsMA7OV5NOolF5ucihWWScd+n+pTNSN+P3k/6q+eWX3bpI
nhF90rxg01q9K3iUFlKjZ/tXsZ2+GYWNe3bkXZkGTM7/GCrwPerFwsU93gr0xdao
jNg4GgctUxYvkZF0SD7D7bhpWHXOvzFXo0gu2aBoUdWfPGVljwn/lYiI5axrMs3c
mGFCWpRGR04V1cuO7LxAS57+rLZ49W9c3UfnXrUii6DcJZKGWopgmo2PpKR6eSXl
rJajKbj6MUVcShCqYvQzyEqLjwdDeZyQthe1/p6xf41VJkr0xhNhn9BeyXbHYu0A
3TQMnfXymdMRWQUzrg+6NOck7UJ08SQFjGM24reTqDMx/jg8zmT/GXCjGaatQyy0
9gIGxVROT2h9udKbB/Wu1tkVmCelzDDSHoi134ecsrSyBCtMnEwLtKHtKwOCAWxS
awyXQLgXKw9EBjCA39cjzj8X1gYcympcX0OG+GpaJW6EPuQOF696omCuUWkslj3/
OdFfRsD18FWA8SbCZOO+13U0PV1SkRe5AXSSsa8j6Gp7kWEEzYBcDZY8YII5C7E7
hodOl2Gh2KzPcN444/aWOsJDOsMx81gy1sZ3glBBpbwAymX2u94phN3FKyFPePDU
ykLFO2ihI9G8Y7dIiuYyCeyE7+I9QRYDNJ71TqYawloKmH/NAKqfzlqBH/1mPMlt
zBtfmcCxC4Z662A8v0o+WV92obLKCHNQb7jHD0MWzfp+JPkJ/ZzYusPy9Zuxsna2
EX7R1IASJBsW851PEbPxKg7gmjMpQ5aZevnzSBAD8Ent+61Kazujmp0NluIjGYbm
uGN5P9dkXqz0HCjymDWE/SF7+r85JjSiX+FSErsRHSjT/vYIxiObCZ8a0gXTaORp
V2jdOCFZlAVWFryC52HcEkBlT2arButQajNVyeS0V6e9HWRSaQvOisO0CH/Z8yIs
v1I5yrJMb6AiMfUNQ/4wbyLjIZbDPpAi98v0KHGd46zYT7/PgiIERck3AJeghEf6
McCPd7WW5pWdUO0dWT6sgOBWZbEXnSaWuBhlcrj9A+I91hW8TPd49Ygdp3sL3jgF
PkUI5+aNgOqFHpx/nZme4isSSSgqaXBIm19wELFF61/oBr2iYtHgrKlGFW+S2+DM
autXgupvRpOOeipj2v+qapJLeFqMAXV5EF7tu+GYogBjU3Z7LMdkC8s2+a1Iw3en
SReEGcak3Hxx6+WKvCvdF2Z7jgVW8DfxR/6G4dzrJ6iSAA3gpJJfORGqVB3EEfSL
YlNw5pRePguURT9w0PBozPu0l9r0PPjD/jGXQmCulRz0T9GVRi8BWTdMZoirSw3J
BLcMOJXnxvjk//6hpy7TDTffVy0x7+sezfwGYS4BdoXZL6q8mAA6xuc3oJMcb6S7
alVg3lxaPTlSHrbh8yutfrDzxdpwHodoI2mPpfUiW7zwSTYnEr/zqI2a8yswl9Az
NLGRVEDfupi+UX+UXSJDix/dw9tfUgCHFlnQmT9b0+O+XFW+pUrzIgnsg0M70RxI
VJr3Uawo5aKzTBK9HeG7MyrOvd491FYHstDOyDHEvoVqBgt3UO/ni/gcHuxpwZoO
Kt45JkoKrZ7Z8WRc/VNDc0sQpS9Rhy3z151cECPeqTqKY0MuGwjCyc9PMs1vHdL5
hqRJauAqr2xIFKCPRVwiE/S2t+HbQmeKRcM8xwC4tfRtsIrnVvWN9jirgQA0PrPW
e2JAwfDJXjhKJkfeIJKtBDVSYSq8OMwRf71y+QDpWmyRBMILse4MDsItnAU1E9p8
5bxl2GI8o1Avrvr+oLBGFswu9DLMKACP0VYyIs8qz7FDEIjprFE89/x2WBeIlMo9
5iW7gpfHVGYx+MgDJdUfPBnAj4VswTQ7FxtFx2IRA8lu05ueVpFUabgGVdK0ghAJ
8bJ4RgvqWCUgvqo1G2qBGZa2kBgZEds7+DaZy8BzFZI9lO1Tf1ftWfDsTS+q4AFH
w7ee76p/sWo4pYuFqnq/gbKh4bKCiuXbNb0q+t3wJ7v7gjwSGY5X+8SF86+nRlTU
/ZkMIMUHkO7EQyAFOw52efzOb8vUok72I7LruCcy0sRcXHPZG9vKiSh+BofXqzQD
nae6OPrD2mN3mBzosudiSGfAhi9AjGqPvnQ8IzvyZVxadKoTOpriTrSDe7a50Pis
PqxN0fwuafUz/Sd9ixunE4Zah8HOPOyrv0OpeqXGgukKlm3KFO0zvmT23phcrYt0
RebSXHpeQHmx/6mbYwwHI2la6CxCGTwC+HBboxlTmPpWYRtRagyhJVllt5HQqIXp
1+5vNup9zCxGMASzHob+MqU7+pohxR6Pshyd9SXS4Ayk4OR8dmlq+HV45gQ/THpK
EcmqXerW8yDy/IHEfIyxxr18qHJrfxd+Hy9WhVlFgDa9gUSUvyR9IWnG7U6eCA1X
jvONZhFhVk27UBP1AAnlF/GzwWxdQrJs3mQC8TwTYGq90kjZCwpmerC8YkJXnRHE
W/CbvDsB6KBl5CBQB8RgBr/vSWjVbCVRU9y5pjpyyHzRN9SZIckBu4GjuK74gL7C
ku631SqM2nFckKnSNZ7PSAN4HGWu2dRKSDm4G2nlSHHiyWlek+qblcwcoKKrbphr
zcwWPZbSVfH3qoGiWHCSjGRJpMhuY5NTGYesuisejQlYn4AUUYdqaobbqizNhziy
VKz9gc+YgYJhj6oFAVhI2ZrdPYtuSUJDxzYmagyvd3YMAtoIvVr963sQ+0Nlujbd
lSy0TPApY/ysqHonMwVpXprSFP9Bi0SyDYD8jkmqV26pSPLmJR7EcENC1wmFdGWO
WoX+MtFcFz1OB6QFzy0tSIM/8yB329tJ0Tyj2P85h7OYPSLRPkLNjsvU8Z3zZJhy
Qt56uACvE3MWe9nxvUaO9cABqamvPjveGjIAXKNL8gFQTYvU4PmZaQ/DWeDUqtkM
wcdRItADmDU0Q2eWQOkDVIswu9uwigtXtXz7gq1hUalsVYeJdUVk0XpcKOrUKufj
jxFGTKBOCTDD5puGZt8cBfbVs/r67DpHc9FcBUxvGU1/BKkLAqqyViaH2gCg1VwY
myzXIwm9y2OIgrWgL4I+7lFLHJ78YycCnyt3J49xSmCOrED6rVRD26aZvclpeSMr
+SYrcAtqyFu5z/ElDeGD7uJLtIIzmhnBOi6Mw2mzCoKkTEkBRoOOwjogcP+OK2e4
kgXC8qDOIoJTVSCYEYUQtfW3lmXsP+6XNe2k4uiM7ksaXkJKKeXG70fgjEz9/K6d
BjU3e+EOUcWVE6a9OvsZ/PJfkWn2BVnGR/yHNub7X9C0iHyfO+9mDyD1+qcZoE7d
uI66m8geiKKGXfOZm6SAZYZ0Y/yxRbnSKdumlR3wwU+jnSP30eoaHWZAZ96oMg8O
585hqdfTy1bM2v09vWg33DDcHF7VP1OKdmKa9lOnqRglqKKbP69iWdyrzrMxlKLg
8QR0N+RQuUeQBIM6A3N7EHtTciKwUI5qHO2uSnB3XrK6aze3xdUHjdoiZrz+emXk
V1vwf7FoEISMVcmoApv7Eqri2iTzUxjtRKU6PqXPwPliZwvX2NvCnCEln9M/16tm
durVGfVoI8mCkdga0xngxRuCLN4GiOIHM2DXQJlH5WIstnn+soWlvagPggYrefzV
YzVAl7xND9DVcOZQLdT3iXx1boQhy1d+JB32NPWlunIDlrSTGZ3d/pMPTqu3Heeo
P76N/Fy26/ILOu+sjlnTA93f2B/hFnB6VpTjLqXWKXf7EIkMQvOgt2zNqSdoCoW1
KHzcZPkrSSutyxqZIlgSgF6emsSvUWWph0y30bi12LQTfkGp8ceqvD4xjEpwMacd
BJ75lLaEMR2FRwq5TlMtvvaKeLtkYZN8zR/We6P66eAios8praSmGSG1sGD+SM8p
6plkAAqXKe6hRcagps6VMWplrxlyxjnvsYIMwn+QcGrvo9z4ysTh4wJArhXGVzr6
50YVKuQsoAjwB5ThslFfiAOsrOW6OPqZa9+477qXpp3gnV0E/F/+txrglbL2RUEv
45M54GKl5ZH+Nu2DmQ7zNT7CpUPkuMbv/yMt+SmFPfqtlCYFxNTij+LOZxgokqs3
FWhJppRjnKBt+JOutPpioRnY3l0sLBteScQN4Wsoq8dGEVd/2y7VBhHdSG3stRNG
v1G/rr6c/t3LyYy4sfjQhSQ0WaF0b+PSmsZOlFDR8N2vENO8XLcNwJBONpIk1bwX
gotvyOTtu0i7zCbe/wEYKJa45Q3uwfR/Tu+ZT6F8Djs84xUTxkjdaFqzT7lMbTYI
ksUUErH9VXtTuimNuNUG7gEvPzJ+CFNj6Fb5ZkHT60QIBszTDCqsZGIP6wrNybvE
jJSVEzdYDTpYlpsqAcc3L5Fwsu7OqQSCMFpX9jscFXYp9/JtYBa7IG9RUqVD6iZf
6khkA3gEUrvm21tJ23IqIbm22FM0da9r30tLleVTkMFGFQP72dRWqAL4BKr50tCz
ZihEBaStC/u41bBN4+85ue7PPJ2KqkOG6q+43dPM5/io4sj66wWJFv1JoVp3YS9O
amxh39bav0g2Q0dKxfD5XP1btkWd440Ej6hpu0GnC7fv0xrTTvqvE6Eg1wvAI7vo
RpqCjF5mKhgM7QwhFqpVw0L2T/6IFgOt259dmXJeqZ8QvSUC2fPs3MwxXeJ7mj/n
bZ5kQes/vn6Y5X7JPYy2dQ/dzQMDc1kGr0gnsdmLkAgis6deQeVJlGWB83E/EOdi
GOlt78F2o933XxdD3K8x3OnoP+OWEF3z5bBu/a9dHmdtnmnttcPrzE7GEqooOaPh
HLnJNIiPMJ4lVLWQZEYi4csA0R3l+CieQJLTchPwsVRtLKBmuXGMZFMlJ80WMJiW
92hr+Os4YBzkaaaSIjQU1XT55DZOe7M7Ux/rXjTKOLGIppXd1qhQ31uIkD6SjZo6
Xg4dirFfNXIhlB0Osa9/E1wUItuVNP0UfiBFSiF6GYcWaOw/rS8tImPmVNK/zHLA
aACBGtqMg5QCD7mjVDPyeDPPNPJdrqozLJeaK3WejHGhR+rJW+WWQM/xfXrIH/5T
w2BE2yWqpZgjvm+imPORkayt2mb2t8l73vvmSZG9lVcFMcXm8UkV82dTcloMdfyV
mjrS7OhlG1nbNQFF2JZV1BCvR6kgpHoACuEaeFv0609tkAe+71UvVACn8QG8iY4g
sBpSoGkHT/aayZD808gO5Sw9sls1ff+FPGblC4gJ72WDhmc21fuCu5AKuS7sEtpo
43/BrtbT6/iZvNjs96Hl848Cm5aHRREDcL6EswQX+eR83it+1DRANLOL59M3oKji
fS3nXSnYqUxiOXs0LwRfWWLUFnjDLAaIZuKRgPbPN9gg4Tx5g34s2Fcz/yKQjtU9
XOVBNrKjUs2aLa9ekxBdExSjKKk1ERiAH3p9ONf478VWDrWOKejalt/32MzG/GdF
VvNhw3IKXsoFXOw2xihFxKuYswiHJRHL54Mph03khWxiro5GBvtij+SMgqiEh2w7
hvcmIfg8Qsh108ke/qGJmHWvepAz8Kza+/+LtxnW2atYKIAijQE5hbhcuhzJubud
cAvwb/XZyP8493796WKxHVjuYI9vhb/2zHssQHZNPjW29yQSN2cp72HRuVKmHdlR
EUSjjMXbwwkgwTxnwdFKUyJvckVk7X0En1pD76H80yj+3UzcXH7Ia9kYI2un/U2n
nQbl+T0HHqAiOEaWQbI2CIGvF6WduR9H35fHJkjieuFXmg7pb2O0ZHxImNpcFGDs
OylllM9MJrD832DVUxPyjpCNMQIKjJSJMxX2vIMY/dQaLZGJEh7REv/rYqd7kr2O
IFVFFydx10YPvsGO5zlnfsCq8wzcEiS8LWh7QbMtvSP1K2ku4tNzRpOkx09JXBck
FMJPudy66eOkha1D8KJdD64e5YOvVE2wQ1U+UtlhgYN/97PKTQI4OievrSsD2oCh
c/fkxd1SxLv/UTzT84nqE/IrMR2+LsNT0ZPcd97LcM/Wy9T4uVvttfwiqOViyIVb
hgxzk6sSt8S/3fPCfk2oCoAfF/fmflQKCGCNCD8ZptvU/X3Ju29xhaque5Xvs8jw
c3E7mLhXjlglSINXR6ZiGB21AGfR6NoL0ts1mwwLe+Nu1Z3fo1Z7QtKMLg00X2lO
6vXFoShpheKbBDSNvSIGBC0g3yok145UEznJJKfPqZN/jRk4NeFY9SlxhHIDBE0X
hsmEvziZyr4HWql6bjGQRBGCRNPalXUAw+5du7rbsvQQY2YYVR6Fhp1BNYNCazvc
TSFAYC58ndOvmKuuNkVp2iy+qzqHtvAUvXVxAJCvjpvy4QYq25H1sZWHmv+N7qLF
ihRMrf2Hu8uruaAgc0lgsG7QadAmHhPQRVn6aSxDeGxdT9O1iTnV+KvmrwDGSxQE
9E+aeAw2ZXvUtV7UANSKZtBCQnswiTc8Ac6+6vSxnBzD7H+NNE6IpGnAefxwBEod
fctJC6o5y3HhJTYfx4mcozNsyjTeUAJrc6VEDs0S8hxrd70gUtqzQ36OBqiJ1s6o
73MJvk6VHDqhnmOci8HvnzNI2zB91Ju9YmWOn+gQbnVNvYOOjP7U9rhIajfr8MuA
loqEW3ph70MUq7TxbX9nHjormfDS5oK2zJMMhLARbVkDoVBSvlfBYChEPTO20Efg
fFcQUT2VovKfidthr4L+R4Jaz/Pm3kparNeyRatVM9HNDsFscYjBTJMoiTRlzNAH
Xaoawj1gZFjl+/Vc7Dqj4r5z7vJdyasagU+LEMDiSnTrLDqsYHQGYV4ABa+ymu8M
+J40+TgIMPTgxrOxSMGNMdNgrsE75fbFm4aUSI4IhxB9utM9Q4oSzXuNsA3uC9T/
CR6fozVL17F9y5uCtz2cuhVz0GFELh2BgNzxvh1Ie14iNw775r50+zFEB98sHX/Y
O6g9mocuHVo5kFGTt85xLZKfAnorL0AeUvD28J0Ch3YjBpPC9K2cHM2McmfBjvhZ
NURl9toDPh9CzgjgX2P4wlOaIRg5faKnHBho72UUkQgwAIvwM6lKzMIy9Amthdgf
DJqyzkWG147xeaZTCPicBWu3JCfHmdUA2smvLOr23fnrNgXSwpHKni0Py2XGU5Fr
EgxfTi5Ojkykg5LDkp1U6x3rKN6203CEEi46UBeHm9MWRIT0Sx/fXg3JkjHFHYtw
/1e2rdxAmry8UJWWSRel4IgZoFMXEDK+5mBip4KFZ1djL+cCyqDrSfTv0W7qEURH
VeO0a7qELy4DJeXaHyLIRFDwN+Uj7mnuQiiWCM8VvTPaFpenYRbai6eWKlGNZPTS
/TJOBLlaEP7VWmMC+wr29LAr9w2vieiLMd5zdFerpn16Vyl1whE4oJ2GDTlDbbMj
8JC6ZvJWStHs6/6ogNdvcqgiQ3peLUzBRxqbGo2yo5DeH2QXGb6HUOerFSRemODh
exLH5/8/wPGe/nwPukbQNzKmj39fHkC0JRu1+Kiu3+OQP9/KRUUgAqt59AvyMZmx
tPeUGjHXF2Hi/cZzuVc8AApIMAP0x+dzBqaBcfzlLOvghhJ6sHrR1tQPvYrxurpU
OY0Q5JMy11ofzOcVoFv5p2JHCxSmY5+27QIARit2ioMhjixAlv8wOGsh1ilHuPST
FH/pmg7ICFRAES4nog77ZBl36a7NUMaihGDj+eINZm6Tkrf7YMIPG63UzA6/a5Xz
8k50EW8KjZmsA7/94UPsIpkMj1ZCKFGB/mZMQP15FFAmpUPdn1c69/wDeZ2fqTuF
IqxGW0gs3HRlfTrakF+VLSUXpA1nIMcuKvAsufDjJ7Nk6gryTeY3eTLjzSqCmdtP
v3w0HRhHjWLMzWXFeOlZP02jQXlsP6fdA5VYBQFaEHoEe0Ajn7FswNx6hS2w0zpw
QY7zs191DU8O3M3vQneRDJURY9kbF9yaJKN1ol7C9EYwQGZPnSrzySltLED8t4G+
oiBIzVPmdPlKqyBYse4wZQ5hqcOpHHcEfEc3nNt0XLkOlptpyW911uw7wMRZJjlD
7pBGolBODFmtrTy9hnr5V5JITFhT3KF1F8iT67ZzZECqxAQA5iqiCW+VGN92JJQ5
X0MNnz9wh1t+SeB7Ppws4AknwNkWE7tFk8cu83rvvFF//onIc8MYiGpy9rSWWwje
Si3nuasgOGro2wij/jAWXv41vzdLTAR3ssbbY3FcTTFnkYrSeuGLuEBTfbSWM6Nf
UR3pO87D46PA1oaXyV/19GzemDKyLmpvFZ4eZqTAc/PSidyiN2XtESZv1UjVz71h
pjbDdtmoSehwu39Nx+nSCbkZpd9buxT+bWuKAfcKp4vXcZLa+CsamTbO7OYosS2c
57UxNdttcGDc7E5xrXPBpnReWuBuvQzgcGpu1Xwkzx+meQua9lTjdovN4OTdQYLy
7vrEG7zjBVdp2C2JpkEBqtH7W/VxeDppXSBZ1+8ZKa+rIXgOh6pO27Do6WR4+/dz
weMGUnd9nhX0R6gQM0sqBI6rqyHT9l7KJ3+9uolB+nG1AI3IVFmGzIkgfKiRwKri
dR2HJwBO2r0P3BjxNutmpf2i4tjjAMn9nC5M6nJVJ7qg6JI+2HTgcusKVpr1j54y
bSuQXGHycT32F/WpYT3xBGvPa5va8bXvLV6VAHoU9lTA4PqaYuflPnzsWlmhdJhG
JM1jYb2V6T5Q32JTD5WZOoKMj8r1Ig0t7t0brfavXRam3ImA5PFlhW+CWd0HHg4u
1dQ36kuikixnrDQ0m+6bAh4qoArBEznpaNOi/IWGWka5L+XSE01CskL254lXBEvV
ZrGPlemlDjLAwCKMWl/Sgla1piaKxTrVoEQg6FnuWhw+nirSD234ZSt5wIPOg9Nu
Ztjcx0t8NfMah5ZdhSHJeGLQDm3CFpKKIepQ1aTxXBkpSn46v/2YCjt+lylkffYG
Q7f19RSksgaQCbj5RSpv2Yhp46LiIJavqboZQEvytngluHOnzYnCRtDE2I4FE8Xk
TTkDXqQWHCWpVdS13sVuVDPNmbID55CIt0JdRouk/fFjmlgq7xaAi7DmE+JvC2Jx
1sknCFZXXsn3FdteZ/yNZKxs0Zsc+DGk6/FkkqBDxYXNkUYVMb5k6neWsiYHVmIR
gw5M8+6/kPemhvfIQAZ7X+YicrZH6Nssn7QvIn58l6VTJRr4jkeExXvy3gtUw7Rf
RN29VWVVFHqfoaa+cPDC1ONnWaVMR/hC9vLSim6KRbymxLhLqPoy3tAASZOCag+C
DjmpnyhUbBgNh8COAN773inPSoPKzu/i4M8mH9d3Sn7eHaPO/ci+aVaW8MXCRmO0
uNGDaDJZJ5bfJmYtiSo2Mm7/sXlfJSaFlqZi6WiAUx3EKPaNUItiVOtMuNEbSyy7
OeZvXVZfxKq9IvS+IwmaOKHPT9IfFQd0uB2wtkQAYz4nmoPGs7GzKYOJuTMtwIm/
MK9mXW4NZjkacYmFgNX/YIk7t56mGUPfHCKYs1k91oxgaRMG2ztxCgl9AY7HloFn
MltDnnP3ZPK7j7fJpc7yNGrBHKj8CIHew6sAEiGvKwaivVull1zZ9QbHjzcvl5KW
/2wD1EJdRI0SIT8k7YOD4glNVd+k9zvHDnI3myH7SEgJrlFW4QIAl2dGkGFoaA8g
HDlzbfw2k1uGVkD8DzsQSzTeyGiOICFdKR8Yi3SVz8phqzFpNJ50Cxf30/suFoD+
t0J0t9nGwaEgkJnXOo4Xd2rNOAqt5CVWoayB1aYhXX4D1Ia0Tz1sn46+cO+OnOnv
lQOo+o5Is7CD1GWWnBtAxOeXagpw503cQbYwGDzAxzPUzeh12dmxqvOctrn74H6Q
4Dzzq9Pwf0sgIwJfMHKz5Re6TIjRCUYEzbS+ANI05LpMazxiZg0Z97AAZ7uC9iwd
3j5aHBYjsRGD7DUoMz79wY7TUdcvz7EmKgs4MFYKMalubm/EQiYt03M6hn/md1Jz
Qt7MTu9d0sT1dIiUHFe/pIF/CTedHiY+OsdmiM3r2qcnCJ0esp0WW9lDHSuUJD73
IKZHhnxMoultiW7NZRjwSQ3g6gTEzop3jFo2vIjmqb1VQ1QFtxDjUmhDrERSBHEx
qbTQu6ojY0cHnoPaDhcC2X41ZujZJDxDAkQuluMnJCVU/1xOZCPO2cbTsmuzZn+U
9eqEwZpIFBRB+9K8z2+Hn5Rj9m4hUbiteJcVTDERRVfrVcmf28Ny2eiCKQGoaV44
7KrAajmSApPRhWFmorrtSESGcMnBnnkcjujFXrs13+Z8AWqwySrFtI4do7247ciZ
i+oDlqY63VRc3ZJw5Aig8kViXdeIOCxodF4Ptt6AI2yapfkbU5Qay0bjPw5Rlhzt
yv5hAs5PXNJSM+AYF154HR+dL+78xB/T9rTbK8jRWv1a4acyaeG1HOdJKQxileMa
n2uX0mJpIkD1R58VLW6G8NzD3VkwuWQ6Ur/1DwWz9qAonLkhJL+MqfYOXShYHoq+
TsxX28gdTbERSuwS1+buNbnaQMIcUmbMoMF681+z6Pc1pJvUZPbuZsw8PvVtO/2P
wfNd7eTXOYULMOXnZybxZZlPBLy6amqW1odGn3OIBhYN1+HoWmLUmb8hWVftWwdu
OUMnbgmOFArLu8WGKt7Ok2aDSp38AfOrU9HuHkHNtaaHOHRvanC8yQZU776b40jf
53zvfg3iz4aAe0MO5UfduueBZGlxGNt3RnGb0NAbCeMlfdTHEL6HMAqk4JrIO4B4
DVIDINQ6GRIacxauMc7vTg8xyv5rHqC/T4f7saEbzHX+XYm9C/iOD0rs1hN5ZpIc
E+V3WdLBjyK0AZau4a6NY6V+FStHsRMKjkG7ljE7UC+c3l61EpDutn4/mZILncQL
UkH6PsQccrXWx9X4/Xk/lSdYFbX820HsxnE7z2I/zugiTexmBzu6VtB9bvIp/GCM
4iRvFGNrUU1qH5BnHP0cJLauXq6RHs4ALm3tfaXx6C08Rv6oNPhzQ2A0x1FLI/qj
gOH2AtVLVW7PjXqTPDTd1jNcdMtX5yD0EhYjbHO6ayuhXW3d3BDCjW8HYfeER0IO
Hcbx6LTcMjE8fy97rkx2tXkcIryeSLr7yQ7kBeLd/0n2VrxrqaXqfBausVk1w59y
kJd6oqA5d16lGB/IaguAbaojtouHzk5G7ENAO+GYxJLeQGZ9/sszfGfdtesiUbM8
nzCJiSKbCSfsXhtKqtuy+2QvKSmdKERatGzf6LzryoMApUHTNta8kFdz8qMz/AJI
YOabASIiZZviCcRr/7jbJbYynxk39TGJ5IskikDS14T89OIc0+8bSeKGBxQ7mZZb
DjeOWpQCRiDr3zVsPRca5EWlw1RyMVJ04NhDhBuAGWA0NTMicuxQH09uxLEsqcOZ
Q/wBG3Mwoc/TDWUDFWTpZE+KZAZcbMtOZbIZCfwf9DgI8Jkl5PlsXUM1chGj6fio
h3avz7VSDhfORXdUMDlD0YpJBYyqYKE/Pcym6jGo7QE/ZKjtTBnKzwNsnU7Tg2MO
Z3kEcP5NdB1nbTPEN8z/kH8S+K12evNUWH1PCibisXPrqwYWLOUNiqiXjtlzM9UI
w2Vy0pmyC/o/txJ4/D/NwonLROVJHtbQuskK+HRtY63w4Kd+Qzlujtx0n32cP+wF
SZtyqzP2Tggiuuntg7yAEJt686Rb3frWCejaNyovT9jsiFSFrPAADpxG7+EXKI73
x/FSVLnbUmBmKmAtSkhqvE6PXHsiykWcS2iBCJsnrO4dsr4FMVqpstR/nqXx69OI
DBWBLyKc6ILR8mNVWV8Jm4skCk6a/KQYZyHxlQ4j6IX++vQYi9gRfRGUoXhnSvUM
aecWzUCa0Gb3117Q1MSR+Y/HHd4x0X9Xma+Ye2UR38Rqk5DqM+yyepRk4KBGE9lj
bhlycS/Fa2kL3ZDMnFiIL4yfEFg0LUm0LRjRlJ4lpeqLL2QqaVjji+nkWlPQPw/3
qjT5wC1AmGITO8njdK+JR7xw2KdsUiYRrYvw/Nyidb3gsySXS5bZmZ74wAxT9tAh
BiEWeFTYur17ToWxzNs9BeO6MbSkXtWp4nII8Y4eGYbOs1vh3QbE78bpf/niCWwQ
9b3yZHeAxZ4bNQfMf+FYmqqp1+js1gGSNIoLzulo1sEogHsN0AtkisNMHWS6Kk/2
GNxPBaaOjVy7x+pNUPsbBN2hS6KwmWNV0Ew3jIjLZ6dj6HBpj4KgkAjuIw2S/Ib3
TCLqxonQJ18AQ2zju0nbWNzyNmqSmoM1y+ZGQYMja9lfqJ++siE6q9hqFwHfLBb4
ZaGSUM75QNKAwecjO47pV78k27C4xuS7OIxwy/hbWwKLpFLEwyJlcyfXZyD1N/Z5
P/+VTmBVXjjra4sIdjaP0xZpGCxn+qQVE7zvHfA2+Tnv1kO9GanGZNohRZCLBLfN
VM8rJAfIn1ORNnOPoA+IojpvXkkh0paQjLZlZqsw+2qPM/7yUhhox6Q3oVQyV/Rj
Ld9SXhSyaYmfot42+iXfaX+k4OLC1qa+0H409cnHnH/RK3uItJ9notI0V6FFcTDd
qMfeGVHR5C0K3pNNA7IwaG6zwKarhm1ULVYcXgMOJ1kHFpp5722/RDpTRzz7+9ax
PnBXrrMZqChYBV8qmlm5ENYt0AEpu5RBdytzhh1CDn+VEiZ4dPCE4OMmY/pXxz3z
9tmrMEj9mVYo47u9FHnSIk/FJ1RbyPh5A63WYU8Tmrf3ksCZ5fRyKKLlZwajlvYE
zjEAynI3JllGD/Fep7OyQh3glAfkO8Le8iY6NeGyqQGCiuPwo4UV+VVcsY1D4jzd
/TPs/N0i5KOLWM7plF0U1RG2OV3gDo7TkeaCQGYNaPrLMiZxXMjNys1ZJ5yt8sF6
Ep0zaSnux8y2fgF8v/kC3LULIZ+qTlvMxNXY4IdLUgQgFeN2KfVrOCs6Xo03cnoP
JA02yNsfRE0erEq9qAgjuCJZkM4LzTxl7zoTozUm6Nu8xQNG6u+8WQgd/BKCv3q8
b+AonOW9I/wCZxU+Rkv9LfZf385r8n7ikl50y4RnJPiuHxtCAB1TM5pv1yCVcfCe
Gjp3FMLVxyBI1hEHZWeCxjXP1kWMJPd7hyCwgWHsXDf45QihjcnmVpbvNzHwty+E
nyGXloKphXNymQQ5xcqGDzux89ACYvZfpTGR3PxLS/cDkDkCNk53iGC5BWxIIjLc
PeSzclknRz2vNvFkW3lgGZZuweDnYk9sCvshoYhvCIiG0Y308q9ZjmVnknorz5xs
r7mxsI10zN4p5aBYkMAJmzDLmayLmUiwGmgzbdn631POND27Ebx0gHA5B2V70qpE
FDJHRaUSLHAfXXkZ2UZFn9F5+lOrW+9dWPG75rsgtW304nzdzE+2mVvytLpZIVG5
40fN9A1p4psWtWNCZc1qYqIkpGTsfDZtJRN/F74N/OW7YxhO1tvs6Ij/s40X7u8O
V4RDoqt+dKCSkZEPoJCGYJ6b25MO9KuGBx+SVMxnDqQmS/1vdtcuDW/vjAyVSa/B
dcAWsHW3Djn95hXlsZgdHq049BnOGPfW1Ap4OuP0nW67PyM2A6o8N94xE+4NjVVC
bMYT8yTNCCeig4rE3dskY3nlbjS3jdlPlWB+n6uG0jxWPrMomf/SXpw8sbLJBFKl
TUBdoeQRM8xGoGDEIMwJLvAhYpb2VILIjbI1fPMl3TPl8dArUFT6PfY7ucK3zvMb
jbHvC2KytAJa5WZ/KTUydc3lR7czvx/Q8Imv7qCx57Kvyn/MBtUEpeZDj2cYd4a4
vYbyetDongZHJnU6dzmmCr4k5sQwxj3SX9bAmc0chsRudJL3S0MhRsvzU/IU53u1
byha8QLUnVsT6wlPIyNJ36o+2SXsKbPC8nwfL7Ms2tqHNcjiOBMqTVhX4swddADj
jIq9ieatEOshuyWU6Xf2enqPXum5FEldk/oRpQwY4F/pO+qic2wiE6rv5wMoBakC
DJtAzLm4OcwR7yVm7d1xlbb3QjLOCeVoxBQoTtNcBVXtHOdb7XQpiRkhq32sOcBh
KV7DZFP66yZOx1MeYO7HMb8rL3Ia6gJPQ/7Oh1HWLGUwWX+On9LYAsZ54lc57Ud9
iwYB/YmY9cKB2Wj/Jghn3dlgW9ecVdwYVGuEmltU8OBPjSO/v6hGTrNJVLbfe+EY
KKsq0pGSaGLXADrnafqrOaCE1i9mL30pN+aFZdUp0poc3EM0QsgT8Sa3Uh63Ojaj
9ro+GNBJBJegyHR6c7JknOBIVfRaD1NTRebQIrHu68sckVMAjolCy7Vw4AJNpRDV
scmyfKpABqxmFjpXZDfjvcA4KMD8vcQ4U0y4m7V2ctC0RR4MFxBOjzWnvIdq38wU
VaOd5W/9qZNUaOM7nMhDCExRbHGpescLH5uHXK0y/8MZwPLxBTA9kDUUL4MO/gGu
ipt6QwSV5lcDVQxAhkeMPB9foRiH+KB0ILdVOVwEqe/aYBFR5WUYsjrJFZc5w2p4
v3t3+JW9ghV5VMmeVLRkghmINgRolGmAerqGUxSJgRT2ZuF136l9iMKndeiQ2XIz
MSd0OTIgu0STy8NXzCaU2RBrsocPTraKHCO6FjW2ESihH68qqxlZQzoAwrjX/uIq
DFqqlDPFK74M0WU4Tkj9E1DSOUAReveKoopojvi74koXk6agZcgIDxvP8ty4unMv
YOS9NddabLVHZelWKQPlWhjf+r7955q1B8O17zwdmq+MTqEHrPf6HPotTTVq0nZy
m+WKfLRtQk/Ysc0C3DrvqLNVDmcs3fGJxOxjHdx9byC45tM8gST37fi47OPtOeCu
sdNBOu/rGzE1ueSDGiHTAW6JpJxcTWxDGuIpwfKqMJcBDkExkVmyToO4wLa6MI8G
J3a7B4/tCNdnn843bR/GnV69+1YL2YMnxYyE/x/NoCnSq/xuRQmX7gGteAu1jURu
Omj3ae0P9/pDiWqkJPFqr+DqhHJW4gN/yIU9HO4gY8/UITXF01pKPzUVOmp4uDvi
tmDP6sRUvn2KO10Bzq1G+/r8DC0kUFWdKsdtUe9Yf5GWzlCyLXzbIzWKPxT483L+
ipdWSThaL/DHb7O3Z9+pKHKg+zg5TvXxBVHAaW7mYJnvYVZ94oR3XOLhRH0O4Lta
TkWGqWlK6nnDH1ItgTmAw41hf5dLmmcLMlpWtqVvxBsv3Mh1D0aIHfxefHXu1zMp
BhZOE1tSqsXuSlsZMzqW/zFaEtGu2dlH4PxPF+o8Uqz66SYMdVJ/hmKSNZcw7bJP
zp3kNJwkHWOvIwhkVdkawGr7L7FjHC6gnASBa7WURbD5x+FEu8VzML0wB7iOUbe8
hAlVRiWXw+QLn+zM0OXiBLpDFiYjdsMau9JY1xkkcFZXwoS51NbswSkwBlH8BJ39
HFhUYncSicHcCxCYnVF2IiH5tXUlHKRQp49+gZ9WYN+2i8l+exN0Cf4P1t3npGVo
mGmQOndjFv/4oR97JSul7CFOtdSv4ruuqOlr3B3EAzaod7Nu44jqM4rfZkjOqt+A
HOoRV3A2o33Hmi2IuGBpyWt+KY4f2l8cnOUNFXrK6vAmdTJqPIt5fbS1h8q7x196
FQxXStd0l7d7KEKWYdiXpOfYfSWqJXjc4smtfRuFePbynTScHQgADlcctJvtxpQq
AIKY8e3FblmTJHAXnUe72cHkL2DrjFCr40o8+Sglm3PKuDDJKR5v7e4nK3VyrdAV
7mD3JJ87zKuom6pK+MZKnEDMfmSLjNWcMOb6LSbKRNl1mXHbWEdDdmlCEaJ13sjL
BUP2dS+yNuViGpa2JqickX8KA2ZifFZHx2L3bXInfzz3OsK9Yf9E/1Ar/IKQcmCP
8u252UeHh7z9gtdwyw7VVY061SyBzH+3Dyr4XHAjFhO12/HG8ihzhqV36vOj3KeB
VWMKNp1mJ44ZRZxoeeERFi8Z/o8VYikdXSxvv0XmFg32V4BOd/41xsGv9x9Q5k3Q
VkCIkwW75a1+EHFsiqUZTLRfQKuv9NlFqsP3QLx7f4gNiMtAxXr525meY5KlS3gM
mr+P+JBpZYNw7QGy+KJTRC3EJ09Y1GGLUakNilsmDsD5VAVnwpZ+rpUMzKSkIRRk
L3IG5MBUDBdrQrz9+3CL6JhCuN9NwFxxWO5JM2uMxXx0NYrOYKktKwWjcNWLYQJD
miutBtN+MifcMJ1A8NnM+9Ia/HITpLudT/Jz+am1yBl3vvFdCiDKT8iqAQuoeZOP
nL61jrUITDkucSAMQasUITdGH3pwlsI7EEuJRZ4aWOppQkpQekZswVTJpu7PBcI+
IywqGHIr+N2ysAPKsnGGSR2+zfcR9zV0Dlgf+tCvbXus5JfvrP7iR/M8nzFkOKWq
JPjl08bz85El9Jy8Kp2NXOroGLx8WLzNJKooHeGC3w1REyBA0ckQ8NhYxfx3jVZU
6DoCrRY+0rnbkkwx/i6FjObkVzQmRMoQfgPlQxeqTBHuj0YrXqjWX8cTEbNR8nuf
KOEg+rNyls8bXYSg8S4ZbKqlRGls1cQVYyMPKXNlDIZJBljW7ewGlNJrV9zW1VGG
nlyHkoEI4YBUT1NTYi5baHC+o64D9sOpRcFH8TtajPEFXG2cARc/+RX3f97CHlcS
9ahV4sTxQgAxGDD7BHTwQ1RALXxORvVhynsrwGLr0XdgD2qR0qfYIZdCM50QZOm4
Fw+4CFzA5gLTDaHckZT+2ZQF4+oagRUncXxEkKI/keQIOzG8u4MhtYh+nVMPh7ic
BApQMfd8WK4y+fLVnr53mH34HR6fyiJp5CFuKBCw3bX+kx2wjgerCgtIdd36YAtc
hK6+LkhgVU1kbFIyrO5S73VAb18/g2GViIGnJ3grLdKP7qjloCM2iZ42ZjBoj/dq
aqPAMZ1Ux3ptKx0qGAxXPws+UeKbi6KHHPWkdrny/J+B8ddZerbNBPifBc3xAgqU
OShuQ/ZNfk0kVqG7nFBNRLWz8eFlfGhtGNDSOsDjP8PpcZ00mr22NyfXk+Hnz18H
fh8pj6pkictmaz8O4riMDz4jYBiqHy/Y0QNhgPFP+rcyzxudo/I1jR9VER4okiJU
DAeBA9uiouf7pK99KQQQUdrrmaKm2ktJZayNwGpLIeFZ0X1BcAUn/ZRLljJr2615
9wOxYpB10UGIPDaoRlAhl7zbf14w0RB+XWb8Eu+4zoqxQDDj9Biy5TM5ewyWACnt
R+K0kqwa2GFWmMGJRJmOWhIkC+84wrIWyZrTt2PvjnxW1C8+KFeEHd4Co1guyVrF
cY3gIKxk6xiOB1MJK7LCcgSFeYjSvrwIhOuAvXk+U8YQonLeKhgHTXpgw6H+OeA2
rMdg4eZlIcuuXiPmyO1vpGmedAv4sfbedQundW6ZXRbtq5lGdZqzZeonXIS2osBd
XpfrZrTPs8m6XzdHeU7pI38bCFdQvytzzKc0m8X76mgAy5HFXrN07PWPlj/q+6p9
XpoqQJvMjjdkvIMewqIFKYPXqVSAFIYHziRMHt43D+P7e1km3kj30sMLCGXKjJ68
W8A2/S58H5LqBqLNMWk5DinEL/niSeC7Ond70sWeT4UmDsf/PN8FoqrO//2QmAuV
2V5Tik1bKo9hbx63xhWBejuZpaoKGE/yv61hkiIJDdMyfJtzNbdz8tayNBLEkysQ
fWuC3IjoTPj93QAdNdgjoE3FV154cktP6q7OpNZkaGCzvUaKomN2wECx4P8pW+cl
EPIrIFatMf9zI0Mian4lWIqGEf9RXV1sZZJCdCf+TgWXrRxqscBiTdMCzhqTzZOv
6Kh5GVYkGZbn56UIFJg7P90CNmpd3oPd4It+lNCFeHmPooOdjcE5ocmmDO8pN1yI
obiSHvWN6wSHv0JWiZ40jbsLYRe3U//bcybX4BvLHuaHAziuqjn3FxlJDyar1pd2
FsmJj51ceDoI2DaEYFd0rMa/c95moBukJ8B7/6ogPlUi4mb7rw7YVVw46LjUKRjl
dSSrZIQhBI7r4svxiJJlcIpHFaBd5+rHGgSMGUodBXHfP4+1wdWruboITgT78h2p
j5/YJ9mj+5qqu0R2HBS6ZL7k0ned8rOeDBE18p+IF7VzRyC9drwmeAkVUL5/Xbx0
qSWl7C6G3y/xMm+pMGrDK7fjpzH0qR8Foqqa4mwqqXMms2CRylguRms4pMvi5/kC
2Z4I0FMbv35n6/IuudMHuJO1pp7oj8coyJOKtoRo2iCPjHB1OK/+I5KgHcVDZ4ZH
qlAbvP/nZl8snoc2DlH0pYBS5N5ytEVj6HxcTPKS4U3jJ1W5OvRGYvRZZKM6rthM
JjtY3l3Ik34o1Qo6xXKnmBotEZnDObMfG8fWCAkamgjwLjjsI1ZbE+TR1XzoECt/
PVJFp2MJx/2PbV+Em9AHSFVZkHG5cxcpnmgF+mwkcNrCcnqpCKcNxXZpPwo7S0iX
SFFFDfMvRbxJyvvfxoCpREbP4Az0zAmmPakXE+yyzAvdDsW7DtUwmsaAmNz2CY0x
5u4cJ7wgCb2gTOG3kw2KLYtEg/50i7Z/LADWpI050LmNEtTL++9/cbTqLzebkCwV
jrYgLqX5R56NNIMUhx6OBCLCnR1+ZavErdyFJhcfcubwMl6leAv5MAJI4FwP4YKO
lZ0KSZBh76lUBhrzxtSlR/AIAi5GsNVogK4Xnuy4G1o4VW09RobhbF0975nScSz/
2Ewsb8qOnkgheyIvhc6sM+2a5thFQ8mIFDuAbEBlNQ5tvzvqsoidIBw1NIycDKv/
5Fn4Iwcmlnhc4N1crU1yo1LC57JgXUugHziQHDZRtFe1Xq7Zb/zMfnDXmnpn1ETH
Ch5T9ldp1H5PLkqHpnyKGzJ+rl1Crx/0rXwAg1/c4KGIUvbLwUvwlaNHjkL9T37Q
Yg1DyIPQIMK3kv6GjjInpDa8mstiELe74wAbZdSIcIc2KxWXKQCE1lGKHW55ParE
KXbkUxAEAeYG80mQP9xQaSv4jf3jTXMeC2ayX/9V34mRHi3r8991Yy28ZxP0TQBa
+rRIIKPLnzlDfv3fdQgUIbG5WkUW0SrzAVGtxe6FokMkT3RJrrMvhqSsvxdZ4zWQ
UVNtn3nnxv5yUKeSR/Bd54HMG98U7trhg+r4WTvuWncT0J/sxDeB0fbfHaNIUQ3R
2PKh/tSdsrTQTDRXULCOiyXD6TgjrKlXR2Xc7rOzVOq6/i5lJBqWB/Emqgc2JYuh
ItAHFHzFmfyxOFypVOrkD8iUSq2YphOOYJhZFDcma7SPzhHfkmXZkFNybap7iy94
4HB5K2hbbuV70jWC/hPrXewvZH4x0DiFRj9h6spEz7icWuLJNItK94v4vkbAK0Zo
OAlmG5LwMOerCfcXq8+qy9rGxGFeKHbwEHLyTUl57aKxpd8ZudyxuBHWkAQMElXA
0u3fhExm4emffn623kI7wH59WL8Z3AsSOJZS45CtLYSxe9uxDQH0dsvJ1E0OLLWj
O4zvdev/1K1tnwaLnWvF8GH1+GtVG6LCtpKfyOf9EyLoBQcCpjnZ6BDN5Tn+3ivh
gH638XQ/BmNfHitvGnlYioP1GRkBVT22f6X/aIchQWNGyuACJ6n/k3ZEgkB/zHcb
iIYwK4dKNVp+p42wPVif/wwOGXeTPQzXOulRGy+ptAXLgA9US39TVPek+tr1Rmer
yDUpgwgBZAaHnHMNocRaWsJTpaSa3KaYVsVHqPMNFeorxbSeRF9t8ASUglx+o9rJ
/HYSBTgelzoFK6q3zhvpSMLOopAAUD8CJ+qrSj2Bi2eZqre6+Su1uKN3+OU698uU
sJ2w88HzOoOqlFfgOtOzdxuvj4dhRMrLtqjAd4ms2sIg9h6izfF8K0foTrwhEfo0
H22hFLV4rfPP+cNsaPbMPsRC2P/eBYDwb7TEapRYEF89U/RddopI+XpbV5AiHz1V
IZoLHcZIkhTKEaZtAhTGyWThnbodTdEnp/ko64qPihaxyd+nfTwS45KNwMDvYhoE
zB9AP1xXd4CTAeoN9aZjkoLGFIYMCvItoOIJFHYl8M6NoVN/J4g3ylyFG3rAJqO8
o03f03ao7edaIvt1D74sIEYv2/zhNlaj5K2gKhxg0tMqi6cKYlQIeS4GzCTGO0tF
154ZjlydLoEfg+cU4n9Xmz6YNU/XwKPdjDuW7TSvzlkj4BuPkU/0uIY6pR//01wu
dOqoKIZ+/K/fgvsSWjoNQrWfCAXCfz9p0KQOnimNGKXiZUBYrwz0mnRCvjQ2GmWv
36ZZpmBtY8BRKiybhnN2HbLukT/xW+3PyG1XRV6MRb9wK7Z1bT/tqW/dKlTGRlkg
2DDcjZQCdIXJeDm1nst5x44xkPa9FdfXixKIdtVo7IFxhkPW7yUvWAMfgSug6BBO
JzHw0h+cdDtE9mCYC1UqaXjW0tyFr+5eeGpQqlWk9HQmOgLYIiHgxvOoQf5U8O9N
l94c2BYc8BDFBnPOo8l1lS7ofxnj3Wsi2TzWfafFuxSROq+fPqK3RwgCC93x9HUG
mMxDek281FjLHjM6pJruFNx7IQBjWCdm60tbyzaoKf8sma8yBKNg3gyoUEYgSh1g
llMLY3hsYgsRNHxAcOCDUZUFWeVIeUFAU7skaiv9Oc0zWIPvFDH+G253cblemQru
Y1aOa6yb4PVOd51LVmJmFrhETpG/7tM9wT5/bnxjQG8RGm2ILWoAUJiE5Q7pfK2G
Ud1SRh+Jwv8OEx5jywIe9BU3G6PvAgOEXaIy5Prl0D7RYPAy8rZ9dr87lcXxqx9S
qJEkIN59XKI91QCawZISJjqfxe37nUF4bH6MiADtzR8UYCtBdcplduynLlLfBYIs
o0m2KM2j5aOEH955wnNdgchyEZ3ma6mabEzrtKWuGSCws09ho3K2vLpIG+RJJPLo
+mnCifUx8n7ELdDxL3Wzb4GF0tsNQ6UUcT3J5gb7FtlPlRbDB3/afQOguQnOzLlf
z9Kxe5FlIVbYJaD9nHFmxqF8Jst2dF+xirjczSlmmvkdp54kdGzEQukEgcv7YeNS
82aUX9p6XNvjfLbacCPcpPdBEi8VH8UrE6aexX4v9QBlfCFbOAd9DckjCcmp+vjZ
oDI2PeeWg4x05YoSUqfqudMXthMnKWkyX6ed/2VkLQZ1j9MWSdbsFHEHfyvShVOy
c4ven12lW1VAIxfx/cNLDTs1byQ9hlvfac/2agpmhE/vq9MMYeNjZVxY2j/bu2lR
vTwKfiD3biYJRCOrmlN6bi3D2cSdL6NTutg+/qUxf4e4zMtmX7AXBG1pQmb6rN0I
DqnbTgZAjdqJjM+qg70s323vIKZM9n4M6iHkQ8D9JoxTkUjWK6swY8P0J3zlSq1U
k65ZI/LDY2F+o9WWMei8j8Ty8XEvZfXFSuV0/AilFswrxO6omJEGOiHb35888KtX
qNQPaBBpBwD5VNX4PVpC8+Qfa8KmMxbwj3LCV4uP0ym4MPGLEFoTevOBI2UyN1lp
Rkub8dtgU8jAfld2/dAshW4W0lEuenXi2Hn7WCmzgNOUUlIRESG5bVR6cTaGt2cB
CBVt4DRE+krXommE4q0KsJHEmVfQVnMgLGa75BfTjppoKRwagZwtDwlmQ3d7X0RN
cyTM/3ltC4waQuGyiOV1UiNZr3M/YHZ29YoZbhwuJegUuK7KGWLNlNzGV90A6AbY
gO2xUs+HXAv6lwm5ufcJXrYUDJuBBs1j+bEuo50XySqn+S/xbbiPB0eNO4psECWm
LQVszTZ/8KfhZboIiDPKmq2HBnYlyWVRoG1WPvQHUpybVE2PlOc/td9BaCU2jO9Y
9itnZn3nS3NzEG7x7W2YbXP7X0F8My9Z9BcUWPRxzVr0R5e2ULlvaq197h9LEASQ
8huFVYMCfYIcl18fN1ZCy6m1jEiBQkQv39C+qQ/o8Ng/DKbxXztIqqOnrU9sByxr
7C+mxTmzPoffr3CUJOOJAP9Jba/D9+Y9b+/+nCWLFqemHbvJ6dN199tw9dpu56pO
U55E3GVYSniyjXIcBaLeYpmSw3Ue3ZvUNgyyJu/9E6axxuf14yUG2LZ1UGcA0PS4
X0QgR+KYXn3+vTpAU6WrI0TWtcmIHtZac0sw3byV553KuMbiT2i1U/k7FT7zY43M
vt/+48dI9YbbyNI6pqv9npy3q6/gPINR3O95roCUcsGYS0sJBl5PMcS7NvhQbrs4
TQ+UC06VFJk0fPopTEoyPtW8sdBYPSQEJpcvPyQp8vKRV3+SlE6pISj9mJ6PBwga
yKd5L9CHU9ZBadlXXa57z99nUuo8vHi9yk80QxAdCjppDF0UEmbrczWEAR6/C9/J
bkE85UrZL7igPPsuI+jZ9SBPWSjAwZNGfBEH5527qzC934dYWkMgG+DHlcIstL1P
h9fhE/i020JH+4NPBk6irPxoRazMrWpAjSUGk3U/nnv3tcZGuxpvv1PC8884xrhE
cKFrJ6L7Zr73PbD3huBemEeY6lXTtQNMX/gSJ63+hmatEilezoMzhPEIksJ3Ocrv
c9v9fKg5DL6YnQeVIR2S874m8r2qC292aiL2JUIMsny2nyPDcuqGdELPnEDb1cXe
a7sfEt4iyVfLnP7bdQp79B1svD1y6wHwgYhjqz7njsAuh1YihM/Gqh5yFPInKbmV
dtQwvmwGKi69DQCpEktIpvf5O3cfqCbj+RKBDMVi/5pXh6HWqsRRJKVq0zZ5RsHP
LnFsRuBm3C2G7T+HBf3ppNdOaYFtNt+kpHYkchB68/ZfN/A4I7nJT/jRaIsOyqW0
pWmwlOCsH5X18fpTUnbOR3FH1YHkV/fD7sOIrzggYLL5hz5PWCb2f2rWGCZ402+G
M1wi9X9Q78McWh+ckx+VnPLPrcFROT5KkEkrmNomH2hwWXVqBQi8b8wwettr+NXa
BkXc9dp4L5ePyNGo4uQU2Tlm3sh/xVIbYr5VLL1ATH8MI9RkpGBAQzy2hY3IE/5s
k54IbJIAmyttTO/8E8MTnyMKXq+Q9STJNF45FrHEzJ0N4voMmPENWq4CxJJ26z3D
nadqqwkJsyiRyuPeXJZJiiSqr/c5RL4pX8aBXEnx6k5Wlmh81NvArIHV+nzEFgV2
vrOnetBGbvXP/4MwAZPI/KwP+PZjgfIv3awV7UNYdTsTzaJ8GcTNfAih1MPGpZnI
FjH1WE96Mj3b2MxzCLJXY4Aaa8xQ8rdqJBqEN9338/8FH9PUeu+UndUrbaqLs/5y
MwnkgPydBrxz6Vjz4hZEnEd0YvfZx7bPJyhh7rtNilEc6BOZpOVauisJv+8C5eGp
QQ7e4z6UmUa8+jjSxlVYji6J7ajkaFGBhuhtnjusUqOoOPhTLiRgAvOqNt3dJeok
Zsp0ejWJmxTTf+lf5Y14tdDd6d/6AOfDlG67gFKc06ep9a5yUetdQylMj2zYyOX6
e4faHigEzLB3HM+AUpQsN2MN3DpVVO/yIHjrm8hzrD0X2TmqV0LnIM+Kx2Cpdw6K
8y+KdmKCUqaqx0tsJsXY7l3tJhEkBntaYuXHFM5aUjI6tDr2MkU4AFsZOxxWl9m4
Dki9nth619jpsA2vpwyn7VmE2dvFFQIGcldeUtNcUSv+ttYUhVhSxGKQYPreXjle
cgD30TRETdbM1btbR4zSR9hYx7qpSfLQSaAVaYsGVrOnhxK+Q5C7nS+TGDH9YQ3f
MgzPlu7oAZaIurjP16YtLVqIKCQsrbn16Mywqq4KqYYUFO+2a0FghuEtuuGT5+m2
kkKG75fX/CH/nw+gnnvncX1GNxovRtX1AM2iw2KXveItkeRxczsC2/qIKiAxpl8j
e7Lp3cRhNPWr0lR7VNz6UOy1kjdGdufE3KZtuj17aw5y8owArq57TY3Ip3T9wtFW
0XucxxM0BvnUatlyHz53bq9M3pyU4LAv+t0IIKyBnkks83DCkJvMFhFy7WpdV6pl
fVDaAq7nPJJghqdFBrEeerncb0RxoBOLlyTdC1YRvDy8CBJEKBL01q2lO4xY4m8L
TPeHfAgYyED8OOMW3gMBozAPqWuvcYouwNvRsNXaPfKwG0JjXhKzzd40ot7Smj1Z
gy5ENVrw8tjPjHHegjFf3+mthO19a2DCxMrAFrtUVAzbiT4ruc6GmCMeZaON02us
jvDyJ2EKck+sHz5Es3o6ue+vhVxUbCPrjQnwA4yX4uEjnNyWllSm4k/oWdkB4XCF
/WxTQZ4gj4xe0Ds8YzmA0GFwioR8sUsebWnRE2wgiz4v5QLp2k/TPYR6isXc2oBr
r1aINftCxJzh4SiLD2sfG2YnvNvEA2LeuCgOxcShij58/Culp8JrC77WbtsuR9Vr
tn9VmVyQJKs3I9APx+0FADLFpflD5hOB0np5Zr4cbupV0RyxYrx7VALDD7qZSX9J
E8llglcJbMatsCKIftPVoQu2zHFVl+yAgVnKfr6xaAIAqz8JBmBcP3ELn5zbDIYv
ai1sLfkKBhEQ64h2W1HEzCWiVZ6q0GA+Vjyo42w/+bDEhTmGbvpPbU8gvdpkGsMe
Q1k+OQbdhKzjXAsbyJ4VKpHVGRPulA9d2KO4OJmcUUKzI0u+wbsn0IbVbAvxk3jv
+SuQ+Mcor2A6FvxDOCzC7vKGfmmr+2SZp2/NcMEBOMBsH+1Z3TjyZ3v85SOGeajd
45BcqDOgUhBcbHfQftOMM12LcYOjUqucWzzYny+sYxcYm494ixGHZp2/Dd7wXQDx
Y2LpD3Uw9vZXBFWpwmc8ClEnfPRcLd5hvriw6AehL6JaFVbC9Jn/wXRTOqX7gBFC
wqg2yHZFJIOAsNCiS5t9QvTUfjVj/ZwSzLhHAgLfmfVzq30majkif/4jb4Lckgiu
8uq6vcazhpELPT/AhkasW9R0YrbLKdLIi1WKtUqbQQkF/Tm7gZZnOAQ8P4IyJm1w
qzFEbmc/NoinRsNTMaulXL+y8Yv73U8FVBafYhen6tJVI2RhcshiTOSwPlGsrgt5
XUaMe1YgCFWmjMvKS4JEG2TzvXMCW95vgX5TyuJJjNiIME1u+YA3YGrxNmZ5fOe6
qhQ+84dMQoDSiXCYaNfj+us4Epo61WMvBU0Z9Nl5VCu5Pl45hZ8dF+ndCojAD9Ux
gzVxIBN0BWEg2uFud6bnRDjPdFUWS/vi/tQmnTOl7gVaN2CqahhyMZMQcu5bs6Ez
jrDBLELniMIKaLUSB8BxOg3RbnX8fnfKLXZ4rCraxmw0XO1vBzcFuFjsDatnImjn
kHg2DdZ/DqA1qasRu3GP+DLJzw8dHTT1Q3AkYdtYmJWrSKtL7lDfTeUTN3qFdVeR
g0ruhZOjBOJeRrBkRS13em/xKqK9gK9Dp1WYjsdPKOQb2XW1n39hSpW3kIrUV+oa
RhzEzvvu0ViN+5zwlrjw0ltRGddJVioElxuhuJ7PmZS4/Ni+GwNxBEWaWYGJFApS
lodvnQGJK6Yn9jTvyHqapC0dbdfs/alJmP8BBZR3hWpu+JCuaNKr+ijlHr/Z7MqC
Qu3QCjgNhYFl2Uu8+hm8Wfkm1tdyRQOd4y6Sk3kRSLtYE/i6Nvfqcpyef+kpx1a1
6YXPCp6bDwIOGAHD/eroJ1zm4yxEY7pEGNfI4kmmgP/P/nuYP23lPsUZAlx+obQC
IdYxGlfXz3K5pKzm2ltQdzduaPValJbVyoUQGoNZDjSbFWXX2TvQUFiMIoJtSFYn
aVDA4+hYjovoq9qpsbXxbKSktQXll0Tq7+waMQz28+tZ2QlSOGV3msVg65c5ThSk
odRxmaxZblYisZxKq7HWyokwigHN1LYo9xYQiU6cvifwrG6yYoObLGqfu9pJY7vE
zwF3NnrIYQ4U0+7OMFNcvOFou71tkVrZhXI7m7zf8NlQfL4opnv/Us4e4pzUF1o5
v8l2TYaKucdQCWymn4Pb3scYNR3FHKhBdlnjQd9rKgfzdlLuFN4XeRwJSJZtQR+n
WgkT/nRcY6xa2GGAWMdfsNzOqQizsWIIoowjJrx39d4jPNO5OaTw15CyAS4RmJBu
CByJAhs6uQhS81PJiWMHiDBZahr0KQd6gaWWnNFYZnIs6K+ZK5hNItS0PTx2dWVf
Xo7rEIetRRtY+dvbAtQlEXQj1aepDjpNXXqcOoyymFKW3AfTD4aEr9OtLxjMutLE
ZFkLo7NooPX/v5tLUtZWsq5weLb1cYfAeQBGZSwyJ2tM6L6yTwl+93ohb3xFXDZL
5Rg+VMsS7uvn+PCGCFWqFV9j7JPitkHvRja7gGhnABeDUXUwzoAgUycUgsl+l0zA
oLlM2lEdO87lmQsQUu59Isyo6oq2R9L6hJKdBLgywTwAL0Iw63G2FUVJmbCLjLu3
gxZX+DPgDutsSDBpjEdkFUQ6Z8w+pzbwBQn/ILTVORLoQXcMdTyCLPBKkTKJFRiI
QB+vgLQGnOzntr9oRKqyG4xqL8pKfQFq5LMw3LeO/ekQzfzjOjYRbu09cG5M2OrT
bt3WlyixxNunEeL89J0k+qDEOt8IwPpHiCInNxbkTtSmObwip5/egUQGVAz1OmIk
ME4V2+jr+ITDl4gazaSdDgKaBC7ZxVdYhnhmf0pDPf+5hEAnJPP9fKs46W+POEF4
QHRk8pNIX4bIP8W0otgjZPnIOD+o9vulJwxNQvhSsEwHHdBP7OebKWWK0AnxiCJP
rV1l6nZ07vMUbJsRziXaRm46RejEpDfaOxi2n2mvQWApk0TUODt8szvlmDzQ5FbE
3RlNSW2S2folW8yyjUHR4nfnuGrNub4H2KDQm1JqnExVpa7f730hfTX9G+BSRCk2
6f0eFFcRDCtEjWwZDhpdhxE9JggsvamVMWkDV6HsH4KcRA1rFOk58B69ZFggITrC
0EYezhRlYWq5OxYdqv7m2+5thjYVwpWCol3rJhR3j2dXYuaOzFE2m8HNl1MEZBk/
uPBOWj9Ii+gIvs1W/3DHH/TeccM/OtZGowwuzMRoCQdG+3yso460y8dVbFChQHSP
O1iu6XlQpl/kdELE5fEE/edC4VATGBhVXB8GCJwDgMPuAkFtGyhigKRZUbQCFn/H
QHhYeTlzgil8NSEXo2afhe8ro70iBn4fMt5OZbPkAUjg20gFjsrCU7Mt3RSxvQZl
wB5KXFOiv/dxdqnE8f9tMcqHm7+l4+RaXx3gngVGXuHkc7QMFlRvEuRUvOQcvani
4PiJB6aiTcSsd0oeGd4Gdey0dZUNmfQqKvgG8KxeFpPpOnInLulSc36ogEgCDTPp
cG1mEhy0ZdiKksIx8wTVNO/nE1J/lrwoPiMrhq/9dCUo+yI+yLNeKZ/+dZogkfKh
rcR2VrasY6j5WDtyK/wHR4jd2QUonF3FWan9TZtXkgxPpKc/nseQ7AUq3rlE3v3j
FLpD6h8/LyeOWMzAaktYVb4cQILVByOoK0jaqUOf8zhNIJzzYu0hZkSPisATObEL
/Z7ZQqldn5Klzrd6yQsUp79YwBUVVuwpzfQsM9JRvKYIuSOiRlVHi/xpVnT47XX+
7Srpm7/wvnFWqL5/68sYb4Xz5ncTyPlpS9LsnYfYIQCowuyHSU7nYjZmMLLa38Vs
1k/nN7YJ7MJD+D7rSpaR2TUF6TEw8lwCyQp46EiFZq6YOVBUMJKG1T5mq3/9lISG
qILpvTQS/F6s9ChLR6TMWXijlWGkfD9p586cmxO/Ul09TSyBb90aTxzmqdV9Psvf
6gnEJOijeCpmHnQZG/JC9VHH7CkkOjHgO9fVxzmpNOJRMotKDg7WMslhb3tHD3wJ
bJQfNXQ+ZXtJLOu7NCVzPUrwDme7YWrV/foBwsDaDfz2+9YX9I1Xh6oKD2K8YNZx
5uukcLPDYCeihmiTvPRZbhRgY4k9mowCszO5ZuEQEDjzUtX8gntPTNCk7wNo0Npg
Vb8KqAy69C/6cxnEZqlZ07A8WSidKZj2cD44rZGMiJLSRLtfhefw4xGC4GxVU7Kp
CY0yQi2rroL5cegL1ZjLkKZtCtx2Wu1FKqZSTgcv2dRxzWmEzQye3Q5Hpfki0PFz
25WrbF9+lC8zeZ6lZZGlaJJ6z8dZqvAjktn6SAP+YjXeVJXVUSOekO8KhHJaVTPu
7kd9tVbms37jYaCwJFuEbZ2u3+Y+0Y3GzkA1cLj+mnSpgZVOBpskgPGYDGxjiYdy
GNfvtX9d0nTd7nL7j+0jz57Psud7Ne0aI2mRWiYWnvuxk6Yt4pyWlrnHL4V+hitc
uUFolcgukeA/1I7j5l6zmfNa9xAESxYntF9SiP7fEoWrmH1GY2HY+iMa204typ64
0jJg0WR3Id/IvRBbC9axxDgMLn/xnutbZVk2PaNcDdobZKczKJS3odGEs7dnqUx9
efXxv/16L3heIIFwvdVW9sAvXQX0xCtab7wZtq6EffDjuKl90GUAiAx39JH7a7u1
2vFGU+HoYDYBaUUs7FOAy933vLiS2hLVs5ET/qO2a1NdMTyu4Pvtits5L74YCj3X
HJlPFmX2l7UHP54l/147o3ErgbskcDn/LDZM0aL49TNpXl9+aiHR0YnbgNVZJdqi
jy6p+Yl2oiwv9Nw1KutOoaD0C7hZA61GUVSdYQm/lyMOI39cjT0F88jK3bs9TUDz
4Z1DndlboSUr160ag7tmNNM9M+QikNGXUB0cwhEqawKS3VQjys3+hLmww+7WEIq1
Xyx1UKQ/ZU6S64qfqPQy7DMNu4vIUOfrq2SOvqZsEJOi52T99P6w0P4bIiuhpZpa
XrSzdk1ti624ZH5E9eWxAGUElRGZw0/5MbBNp3mjCe3QHrhdD06OlHq+e8LpEW1n
CSUl6T/IX8I31mh8jRr0ZmtuQ8ZhRULdc2mUAAFvaAyJEv4Q/RM7z4/4bSBWks3g
sBXvedYj4zfO/Nibi5nFEKUquEAHabdCGQmzOJ6Tl3/TPX7++ODL7nxli+9SotWS
vnphfaUFTs57lHcgb4KBsY0ZciUC/ZmonT9j5JVz1T5KVEbLxc9ZeeV/aazt3MPS
KvWQ5tkNhBekw0ybm8T6F8eM47AQsypFAub4V/kQSNs4cPQ7KPJ8dMR4z5wOtD3i
IvWHz2dSyz5YWdXqoRcqYGZuDNaR8XQgwBuXgq0/0rJQv9O/tA88VWTVKC/JKI1M
iW4JMocO11e0awMYDEoXqiPEYIjQWb528X3kMQANiC74q6kA8i9HDS1Tf51WvlXd
kgVjrcaGWkXs9rsLYqGrYhatRIScone2wp0O+z65itsINGTlV51RHoKCf7UeJ8+T
3sxzPzSQd/+02mAY7q2n4yPlHZDgn7ojpZJXmBTOB3puGJkj6v57vKM51Av8wDbj
+QFiH9jyHXUepU7qfUzgo4odkjXi8K60CgHxk8Ih+GVX8XTHjE7/5oc67O/8dJ6w
8Z8BFzrplexs9v5UinIVddHg+C7qAFWH2JPFNmNAeEQ0Pj6S1UjOk3fV5zEVEz0o
E/r9kCaZI1/zoYc30ZjyA8hMsJFDOyU5Vef012GcNSyM1MuIJv8llg4UhHzgtuJw
nTkMlDQg317L60gReyl0lHFvzYQOD7B5G0SPsLze1Kgfn7B1fUovCIgY2ysBA42w
cJWRrLjM3bMMgCxsAOTR9wzFpySaPmGT+gXUnZRKMWp3dXhHJMEL9VbdOXkn9IUp
`pragma protect end_protected
