// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:52 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g8lNe23LeB/aOCqEw91bdiOH8mMYcd+nR2Fdw9TN7KmNR8rIzANyayxMZIo9UHK/
91hZQSdmyO9oeD5NewF9NL6HIaau+iE5Mi7woirurAgu2cNGuBYN9bJKR2qlFaed
0D67JChwsASUqk17PJvxNQ2hz8soOsWVL8Kk+E0hcxA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3888)
+F0qfKokF8PDkRCAkzFVjTtVrFMs1vFZGdckQfCEki4ovF9T5BZzc9K0oR1K9AXH
RoBPobPN6roFIFI6nsiQdA7VEZRtNI8QHyXb0WKYJAQZR8R1+1Ns00grfPqTyfMB
4EApMjabbpt8Okjuy20xwBikThz/TYPexR65HbwdfXQGdvkhDGONK8L5JFkzlGLL
sPNgsJpurPfXWdGtrgxsDFrfnMrrCHHPgeY8GWghBWhwH8VcMvu3ohcbxOLWpmIP
o6rWtS5Vi6BcLi4RbConJJu20TVRZ0NpWAap0Al4wtQa6gIt1omvhhwGeKaNiLy/
Kab/cqERxn/aGPCKykP8GDhoOdjWX8RU8V8cC6j90foAViDkZgRpxAeSBvfF6MhM
E+mpz7pfVRP/m0M5YB+/VUEMcq/Yb09f6R7OrSj8h341k6vPvPyELihh30S14BoB
VOOuAZY8v+CajeQAOB5itXfelRlv5Z7O0e6PQs/G8j1iaebfEaF6UKel5YVXbwld
QpAoe9E+YXS+c3L0tmBTO2jPuXTauXIsQNifhMdQz0hBj6GuSmT7a3tIEc7gYRhH
rYxZc0/4p2qeSBEwzYmGo1docXxxAjFFN+NLQOkYHsf+84OVnIkYb3f0Yzypu4Qn
MosXDSHz76CtDDldootEXoAeW4rFZRGJ0fOSF3FaR7LAOwqFWsWPeMZnUtMF+D3C
yjs46wOJN6TUZyK7ISTfWsEE/DhH//FQz6H/ZQwav8LL6KEuzpXgz2/A+SDt4Rqf
/M1b3+CVG5gPxBZmivXmswel4wa5M9ccGu61ezmEU6kWrxTlWhSuiWPQERCzby2B
M8QGFW2DU6BOyws/meqzIC5EnpqNsIYNEJzrtQMHJl/9eBRkifFJRjKd5OsBc8nK
yNjb1hRMVFwC2XH4RnlrhfPhgpIzBqsAGUtKn/xvk8wpq8flM7+ZsC5TgYBxCkcF
cWvWqPWzKyErcU0hP6cKJWWrOnSOlo5bVj6v2R4pQgtG1dGKT6q+yi32vq3mU3n3
zO4S69MIWpxPXGiSiy6o2PoTEjqpuPu1fDasldayX2/ghw93uQjEK0r8JWycwQIF
g5J4qmJ18GuVXjRsdljmW4INawmtPQ2791tiMNZqYWLgkRyA2sq7KUFHjvynhb8C
9tv/caMJuemkebzS2xGWvkBxb7tYziJkssYhzS89uUlQq1BcTEGabZjy7N0dHoHz
qjrpOQSuuKdDUfMyH9J0Sdw0lnG1Jpb4YCliH0euZ2AgKUdfw2+EWvVn+ukonXWi
7HOiL8wnWq1P8Z5RXeiQ+Tg31/VcNCCOUK+DVwUvOEAbDEie2DaaoA9Nz6jlw9ds
wF1EpXqgOTNS0kO5DhmVjkz8BP1wLGNYxo5ly1Dirw/11EoEKjuVck0i7U1yO7dD
P+VmzbISnHImkkgI3PZ7k8aASUsNoC2K+IcMvRGDc6/uLJJCtNcU4aodaJW2317c
Nw9SSkWFLA7weBWnVj5ShCZuU3T6j1Q0VaoG0fZpXVKOydrE0kpM2LsmhVdVX19x
Mo1ctx9X4JkHID4ZCOVRKd13gGfelsZPKH4M17bazUphgzkC70MpSI4If0CWXJG6
ezb2H5fkAAgXYY2AqIYFFls3dhXFL8A+PUXDk5JSnaX92/SAgO8IADxxNfW+VOIX
ScgE+igTksXIcFkjB0AlwJpzPSgUCusIe2E2GuPiFV0gxQ3vsSLdcrUtRwbNZugK
NGG4Kx7eowb2cWFjCRAgaGptan6nAbNexsFyKhKI0sKuppFZKWU5U2K1EFP5hUX4
xacDtGmd7Dw5n0kvY92LJU4OwU3mYSuShFUqpssXo44Oa6aW2IT/z8OV0s2QqZQr
n3kzuIRgsBAFgOvK4Uk/96gBTMnEboEQM7iFUY+5hp75j8oe3+sOKmrjA0Qyeeag
xCsWKnFZ8DOCc/rvyQ+w1mgYe6Vs8C9Tg56HBjtbLuk7lFw7V1sDg8fqmO9bFRY+
3KJV9AHHlDel0oXIJMqcAOd9npPgV1UqAkwzcn6JT5EDi+C3lbyQPpVkhIH8uY2K
71W8lbNOB9y+5sFOFWoYm0jnurXZ9z+aS4Wftc5aXUDAu8CfvLMOxadERRpfTL4e
j+MJgyFbEa6HrukrKkv8m4AJacvMFW6oJxFaFUXM7jX4LRA5RQAVHMs1NhUv4Esn
nJ/xNwJSM7kHaGr0xZjy40ll0nQ1+zkO2UeoQht6j+1GBkli02snIJ0zKkjc6Xhk
QQ5nSc4+CPm9kUzdjtzcs83eOY7hjkiPqCSftyQfSDlBNcBFg5kT8vY3G+6WFZ/q
WoQK8oXFUYbqqc5g6M4fM7T+GjXzFy4yau+vcKqcEe9I6pGb8ukyjoXXisTO5YwA
6oQCOUuwbTlhPVnuHTWgEmagzDKI+e0f0FBp3LkgSqCi4za+yemN3owUP2SmGLNI
vbyTL/7o7ttL9iFBfyvwqzDH0WU69Lrk/nXzdHE//5nosV93ksYvxsKjJk9c/3Kx
4w4nssFKBhKq5u/5s+4/tDS2PjRfC/OLpOAyNg4lqcWC4mGC98D/rVc1p1w+v/O7
R2ro17siaLRnvW73X3bDWBo0V2nw8pUuTkGRr0ZnoAvtmTGIaPJrrgoFRCp/7nA0
9DegZL/lS+SZ8pVCunpHPcB7p8peSm7a6BLU5iaHy08GHiuFLMgVO+TIv1ucxPEV
jg/03SrmE7+yogOPpSUe/s+AoVy1I4n22PE6apg63NnftU/8bksDdYYQuHftqLxb
uQSV+AOS0aPrWE027G5O2o/voU7PWN/junOZlkuishXUAV+jC6UTxzHRTguwQbJt
Uhm3Tf+al8IsUA1J+KHHJiwoyz5GWY8BY/EwUsepVgjdHmkVTaPJpwauAkUbaBxE
jIgTQopzwOSX+fc0OLLSj45YoPx+0gSKfpqPJzKZJNVnMQDfe12ipvEMde2sfxg6
XD3ETi1AYshpHquKbDx09j6WEPfXjRWIRc4a3vsffvBQQS+xOy7/5KK2TEo97y1n
y200YTOH25XClOHISAys+61Oo7C0xb270ZgsfyTKJ4768vqnnAADVpX8ou1dqDf0
n7AHjDskR1eeEdR5E9+SWqfJ35fkicGAJDvR95JwDbL9Vi5R0j+TzO+mLTzLYvb+
tVcu15LI8n/aPheBA6M7nJcvZSamifmFns7kl/ZES0WBAlnLzPkD9HUwZMjgDMQh
4Db9bEbraA6DYU+1vDG7R/cmgFs2xgf+xFTupUx5foKlbPIUy8FUPCjQMNnzbJ8M
kxMq8+2J++sUvcL3hiWIFFxBkJ5bPJ3T4sevNZLtq6WyOPhUA09RS8z21oULMyNs
veDl6Yc41KeEzx28U5LHTCGnExOg97QxwF9BEQ+cJemyYMvQEZihJJbatjyIWNhO
Aa7WpEjjPmDGaPJAKLp20ibSRe6pCwVrPU8HaRnrJISAV/14HVNc++1K2q/VCKzp
v3Y8Zqaxc7qSnj55p9cWA7o5d6gmrUW+lCjVvGkyugNNys+QUkiEZtpKfWt3OkaB
kpYufdeoJspHiZD34ZdrcnN14adtsJ2Fh72kOzffN4e3MvxxUZ45fdbBy5K6qcnu
JsEyonFilZA27LHVOSXGeylLZlpPbC62552xHX0husYj7r86Tvy2+KsevMDgRizK
1XOHx7LCb4UJS5yNrU1DXcv+u52DTSc2im+D8kAUKKVo5vLjv/giGrV1svgvy4j6
I9acUPXYZ4hemYRUSEM/EeoHVRrFQJixlY+oM8ycPz8xNT7YrU+fDLg4/8U6As89
QNQA4ldWnAXjUvrH8AxaQa6Ia5cGevBmv09FiLDFLUwZpTuohIEvKoSv3JGOw2yR
WuNf7dVZ6wx7ztr1erJcLF0O1JrCD04YhIwc+z72+dWCv9BQl5qR9DktNWEmI7Sx
dbCI627JwvbGB4oG+xCjq5rpwqKw+rEYpJJAIjqM9qPwQVlI7lDJtnIXpGmTkGtJ
Dq4Y07ZywDOagVXIg5hLg3w/KO1fZozIikxk8XtcJIK8tCL8s+gMVtu7R8M9F8yn
OKhK1Xv/3WNi1M+wmeKdE1hL7/e+RXBOKPPHi1iSyOv/kyhKjJ/m6QaDGxI7NFwy
rKXGKVKLcFp8wlxPXLMtMsmCEp856Bx517Cx+FwwPgrZioMqAy0QFrOZu7x69SNC
XltEGbHfsJsz1aqZoaKFUm7UqRiZeQWXDJf+5Z5rogZQy43hAw56Yl/azWreXhhp
kiZfdd0a3xA3uMUKnSGL5eMSn2OXVzKJwfPYuP56b+xsUSLKp55uG2A/363DzLhS
CJ54aMheLDVyTITWkUfPZGCzIP7fIqo3aJxlpJaSTQARE269fEqASmnBU5TehHIv
sD3lUH9fOnevDJ8bU/k0VVEqzeuNcVTKEmuWHEPdOjFh6V2R+Ue12PXcBvOiELD1
blpFo9mbTOoo+WAqTxdqG7OaEKClf8P2ukFmw/zlFOocYiKqp7R5Lhb/CZexWVRS
kgoVL2VFft0IvDWKarbvck6iY/0O4svXeZZMu7ZYZdW861WVCsBVK0PxlOO0NOxC
Z1w13NhFnueN9OePTuDRsD+d8bx7EFaMsJpbaaKJxmgcm/i9i1KXAeCnfQl0n+/D
q2FLfUInvwnJp8DpAaCJ6uQRc8JmgBW9TTK7X0HLf5GD5tOTahyTdbAak2SQvmk8
8Zuy/IA8Txb+4QxQW9bwfZ6leZ4uxqy54RwpA1R9FqkZylJEGg8zopxinuRJblfa
G4yHOajGCKRuX8geiMueb+bAK4K1WCQmAx8nhYV+AF3zdiby/hUdINqKKSbRjS1l
9xBsdv87AVkMAasl3GY9gmuoxEzBP/v+veSKefsYJNm7b7BCzpXNT81Zm7OGMaVM
N62myMVAIgYha0ka6Ec4yziJrIQ4pFzcIz8YRijZBbcGpNV6Ms2JM85t9YgruGhk
pJrUJzWI17aCHquUWjmdr92cwysy8fbA9o9bie58LNol0xrmYntX9Vpi1/9Nyu3a
zByRg6uBFdZbPPmvusKNtPsQ5rUfllDMIQYmaaX/M7z9pIWiq4ytJqEDVKambX36
ozQzyKhBVjB/Jh/W/G+F6rhi+JsaxNMH1V9cHrPB+CRRHty1R/CrGcdpfquTRRlI
wh8/uaAvcFKiIVJZo1U3eLE4KyLtboFhA2mVoxPN9jhTBvwwTdesPm5uyM6IqOJe
`pragma protect end_protected
