// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:50 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wd+a7Ud/w0/FUiBBm4O/I6EyzwlqW3Sy3zGS5xeuTwUdViqGCKfx1d4lWjlRjTN/
2d2uQ4vsss4yprJdslaw2f3iNT9DFwyOmWwSb8ma0eE/k8xn13jOFNkKVp/K57x5
6rgjDMu/TdUnaXcZYksWBs1RVH7PFwrM4i1UdUMyh80=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3200)
TrYGt4wQAm9mmGh4w1J/39Ybc6rcU/9WYgNC7TBOaSIVOT9zIfwpNOQb03TaUtQN
J4oL+A9maKWhDOF7XtByHg0T5pDiAZOYbik6wV4GLEW6pzHZAi1Z2mNcZeHj5Un2
KXSdxhAe8i4H3vH6t44hk3rj5pb8Fw4Uci0PKak+8lPoZ36beBWY/aHsTfUxJvTo
bsPwXg07XTCqM/27V0N2IjUmkz/r/KPpKgzn6oKkr6p6l7iS73PudZxTCD9ueYWh
w74iPoChzvHZ3mFcNwHOyHjxIVVcqnn+QW9F3Uld2XtBhw0F/JGekz6/ECT8SDdW
8ioMsyB8U3k6h5PJdpMifCthuEzSV0n2SM8KKz9JogH+6IDpjAuMd+gpCEc44/pk
izZWS4d+wCKib7oEIRd105clTzqUqOvzSPTz77ArTORm/3s2PQqMvwN5CrILH0Dr
P6hGE+/NofCev1DFnP8Ta9op3VSq6CEMUUXmIsv1OmyHLa9rGYD2omj4Mqz06fA2
UU12iE+xNtGrzVXpUCKafu81mPWmgQA+9alO/WIm4g2TnsXbkZ+VMeSCeJKl8FRa
/WMc+EHdFE8QpHjBAz/S7nhNWRpSkh5yXc2wism7GjYUiPSD9eYXxVnT3tdkAAci
MI4EgHTW7vbFp91/vnZr/J3nvr7taBa2/eBiQYuqRoS4ZqNBw+13spyd5Vtfp/G0
OZasEKC9nwvaR6PyeIsX26TbgrphpMYu7qRLOIm6Is2Q4+UGN2apGqkELe2ZBiJJ
Z+OApEqO8aImlfLKLY3lhIk5mC7bLr56wNrIToDS729AzdfjDzXeofdRSdxujUF5
G1D6G2Alj0aaVgWWnNcDKKigWowHsNi5YXfePKEE1Lz7wMd3hLtZPWEvB1JZEQB9
X5hy4taVkRmF3Rb6zUf1ugxlRiVzasxZMViOGUZWLBmCUnYCy9CJeSU9L3zFbXrJ
nFAQTCW8Pl4q6+GEEUMUrFEzpsWKdqg58hcgn6qltZK3hhgsb/Z+VnjE5hnsZQpf
gjeNyRXf6opWGXjdisxcSkuQGJrv6Oueku0KMJL8H+mUl3Kfnm+mqYdA74cfvPSF
S5dxTkBVDHwuAeu5VVIF9kWmA+GQNoobivZq0N0EturNDYDuwyf6/xxIN0ANu5YW
0z9Xk5d+FPVUZjqkl7+ywcx95OMY2NnOLA4dQrxg+atKpscw+zt1vZtG1/jc5U+t
A5tv2rPDfRjkgG0pjhLU3H/6BpGFFps34KAwaJl33yPTSTrtMJpdY910bZMrpstj
fh2POKQKy7Q1vehrYYYheGeiUC2HMC3h7wH052zZgXtrg9KVReVnzgsCQENqvs/Z
6kjx3KHu0k+Jn7ak3cscsdEq4Ek4yIxdrRsGrfpj7AaXNDosgrIv8PZkmw9JF1zF
TVXtE7yay/xlHMZeZvgOd7qqcCwbEnaI+ElJ6JSgVP7CmggTgYnN8CAUaxK1dSfG
gF6F6Jy0uFyXJdIKR4Utgq1FypSNpzgtA5xi0X1A+r6f++B36zc3w06tXYWUYiF5
KPf2YoqL5aSsChyTjHCyVE6fnNmJS0LGMEpkLfTYAonsKcGYAW0AN4GlyZbZeZWu
91K/roln8cN+hiV6my92M2sztPltq0ytvWE3DlbmZRx4UkR4t4yQdmlybW+P+0KC
mCYebyE2wQax9buYtcS2U1cE0yerQlW0OkpjfuAcjD08HmtiEKndK5fpyR7c3I0A
mRarFUGciNvHUqZPQwCKcjnK3jqvRrWy2n51fqY8DaK97Rh3L9SupL0/TiDHLfLF
dZ+LAx5fa8mtb6M+btym+CBpf9oP4oSKI/MEOQGM8y4i5CxglvWKGih1VRQIvnf+
N18IDgE8xEusdp8MnxHhO1IEr5SgoCkb93bX/nyTSlXozEeWVAjIloWsxuDAWkcV
A8ZcV0zfy07gGbEFIJbVTgzh0yOAzqo91h+UMtu5GAIo3lp9sGAL0CiqRWb77tx6
chs3J+1v/m0B5/HAK9rtjvJgwbUxsliX8AaPQ7D9S5FwS3kazH0Yk8CPaH7l8zQ9
aVHYFJ+DQMBMl0J8sejIfM1lsfCc45KBYpOOgIYJFaK/VBbSZcld51TulToKhjNY
MTv4YrE4auBp7HDxWirJM9KHqZa1vT3oFOjmPj0UqS12IiyWnj0ETINirBNfm445
75mC3VHJWJQA6C0ctLW5aSXOu/JCyFS/KLpk94mn5FRIKAzNDHVS5LmBZ6JiSrNr
EPKbnubRa6dFivwLGTzWbGFXDO+MMUhaPo5LSUxyH7W+iCPnMJIfIZ/PItCmCSw4
zn7aGH5HcGCTlW7oEA54ZPsxi5B7m/05DhLZ8fOqH2bO50EPL3G3Jyn+DC1581Vy
6Mz1ChaksKvljm5P3MuJVCESkWIwv4nbXl4RLl3ZwZ8on/mK4H/1xRJCSU3NGPhm
n4AmTnuKkSZm+mdxJJvGeSiDCmjnQwDk3FCVcY8yxlX0YS5uCMZKFJo3qvMf6mG1
AXiAab8PMfjcXdzlEoaCtgp6cwu77z0xtA60NglRpB23dYkEpqyMEBM6p2qsRpgT
FvtV6WGyguRu00e9htvC8ovlOAw+pLN154KIcwSzkk0/bK2OmG9o7WfoGQrJH9c/
HDlF5KwBxm7CDpgIyRA3gtihc2ZjKfxD8xBNmpWBKSnrzyfcv+krbntDuxKt5baa
Yoz9OWC96byoiNjWTOhEHqieev5rdUaTqK2V0UUfLuUVK4yGGfIHnj3krPoWapyZ
/nnCjiH5/T6DmkZqlny2uLK2b49z7nWjIpFVIs9ObSAw+Jx9EeqYMgAe3r3HYv73
6PUYrFKMhuI6hvZyCLxs47uJ4I+eiVvFNl4VRvRf9I4jUysQIOjostXukLuuRtbk
rk/oMyU49QWf+BNFuYgE5jhh8zxaStv0cBmboTE4cNTZx3eYeSWp1qKWGaJb6Qc5
GRn6P5FoWx7jJQXBTaw233//nH1pvU2X517VMa4aWQW922T9xbFLnJshbVgGp366
Weiwz5cfff0w5+I6uIFawRvvHGIkrJk1N7mt1ddrvJAH6DTN1ZFGsKkh6SJE1eWB
5LhQiiNScVDCNHofvLOkWSHR+fGRoFJ+XAL1Sg6sBKTkUimrc7StmbMw2CfulKXn
Tozgw5S7a+SWOu8v/RKgR0CKksutrfqPTDXy80LX91uYBrTzMb7piuSQWb9+QZG8
89mdKxg0iTooVqlWFImC341Ys8ubsd0pbFQ9c8bHMaTV3Nva/gDrE5PanDRTjQqL
ttgm+7RWHGZ+EhV1QYLrUUjWkCHG4J/1UzxngNuofVqsc71WkE1yzJxJdMDErKYb
RtVdfaRaooEOfyzBrvj+t7ccyez/YRI3tIaQ1NXKj40iOrl8edGgzqryzV4UkaDc
kLXExNuc8uJzoAd52zB4gMEki6NjPvgAW/k8CFwC+XEuCG7wlsfl8bf3ae/B23GJ
4xYzA914qrd/Kx6q/V59U4hGXCBsn9YUrnZNhqRMN8yXxxH/wwx9AAwjczOe0c7C
o//G9lqTer6GdfvrYTd7KcXrcuUpwFdeE0JrjPfAK3oyPGAlpxc7+Pvht4ebXFDu
k2+cugwMdVxDuaCpiqZ5pbr8TFKPChKws3vhYGh+GWuuLufQuCZSm83FUCop/7+9
rY2bAnfQF+Syg46URl+MjBaL9De5Vi3As+RTMEhe49eD3GjAOaISDQpWONyB8mPm
KEXqwgbAqZmNzyi/Up6Za3TnRTbPfw54c2Rtz5lItrGcKj8u2ok/NOO+EGUWkSE5
zpDHyhi9FbCGAfXyyIZC/P15KFxUP7WfA6M0ZBJEnphKfLFquprM6oiZFNZusIgq
cdnXQW5bcow7E1khwhF+ptG9jCEleDzA+Z7q5FQ0TiLFUuqR0U8HdUZXTGVcc8CV
viBPC7JWplTSArUh0e3adzxlJnIGVAp/qaGGTtxIcA0jKjlW1cauMiAn9qA0V5FU
/m4nrDqKcz682ZDyorN3cOkYi2O67B4iQeN8ltUCaMrWRdOgp4i8eL4K6KH/2yh9
6n4spEPNl3DlbPPQPMBt3+XdkneEsjdqw7O2RnuDabnqL2USc2QHL9UVPZoqEKIt
zpkhbd2Ti1SM/kVkAZ/P4abFdF9bfOcpHsBov8JHUmDcBt2zQtvxW4V2amcVYXpl
rQOIeEbMvsBkkC8wxRypHx4sg7vGfxK7a1WKypq0/+8bjoLiq33X3E2FKMyxKTMG
VMoiE6Lb0AXnkJ9ePySolIYTBsV3p0uTvG1Ektcbkmo=
`pragma protect end_protected
