// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:54 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iGXj4ZtWl/qwHAvjM8Mh3ljqLB3GpIa2MENQnhKx+Uj+jriBa8cvdHlKrICGusmA
8YKEmiCgcnzrpl9FKzL0A0uELmqEWLdAuAbz+M8JpwKitGGFYsLMw6J1h5Qq9wTe
7NPQObAII6RpwKZmaXCfP7T7Wf2JmGqnCKrg2uf6vXw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
Nd8WxkZs7dLB11FdcojEgfa0SuT6CaTkqRF0L9W1X+XdKweo9lDUet5hWJBxyg/0
1TsEYG+6EEMSecliv1160ilzNAD0MKS63ILxpd5shFLyy/Z64aNysLqggq6nTL6i
c7TpSxEH8QFmLcYDHkHHXuQq9/Gwz9IUf3LotPLnjVkJc546qNv3lzsi6iaRO3kf
9PT3DNqXMbvrT3MJu44XoUUtGotOgabTAq9Wdf242tK6s2hTvAGPMcdIimm3TWQy
uMxWRH/irRM3VawiNyqkcAWirA17bX917l7oF6oS7R4TVCPN0cJ31xiCLaNxZkyU
ZRBMZjed0soRBHDX/Z5BScGzTdwT9YDl644dmqtChhqvbjVsJT75+lFKKrR3X0/U
41RaxR98llV8KyWkk73tmpAaNxIMkIAxMdteCwDJpwQMD8mwOosiqmWZ+uuZVIl8
kaSRmDWj3C1lVe6ioYmD2+zv88y05eBpjk5FPVgV5epKve6oPxnJeBArxFkZhO/g
F7z7iprndXbbGvSjsSOppqoXCXpthxw8FgVikhqkIFk/QFGlLdFBSAfCe2m9zFH6
HgqeD9CueI0Hy65Z4GZe8sEWu40MNslS1UfAwoSKoyVm8n3u3L6gmuCtc0dzBX79
gLgDjGVA5n7GeNK/DRiDGhK1klAcXvYnRxf2jNfwo3S+QPdD+wGLmGIJnK2PZgrJ
fwvPgu01BOekj07XqP153HQFQU0zxURAaryeK8ML6WpX+yBI4FA7dbPYy9XAtWP6
hAq9vA2iD1r502CiDjamAlwYzHdjShOTY1rJURaQvtpMVWf9GQx3XpiOGPXUAPfx
y3nwPjEqQapAeAO2k7Cr68lwp79B15yaMq5wqzYzHQxrloAcXAcP5vK0pf0N+9LR
LzRGvg+IHiFVKlhCuBEi4wlUgEnlBkm9Ndi0FbaJQztMibvQhoukCkJhe7+q9UbJ
eBDjEh8VIhZ7EShplmiqCtvvxYOLVSoMGBSDYIF2L7VwZblJ3Riexrhy2eSlr8L3
zQHz2ujJ6AgchkGog2iCLV64MOSuZY2L4tN6/bWQu8WP3d1PmGVUj9atKJrVs560
/J2HZFYEZLCWW9RiwHqdPeSnmpTLwgx21crrSTpQCm9gEKOYvLyuoT5j6ZfsFkqj
9LbJ3B6+USQx4aGcM4b9H6bVtAocx2n2XsqDHkco0ML5mteSNBMZaA/lf75UqxC9
JSLDMvQMIASY2JWgFKstkoMrs5GHQYuPwJ75/qqLiMcEpOfe2krAidpdgtmti4wJ
SnXtnya3IbJTBQ9FDiYHaU5NSF/WKwPp0WcEhxOm6ZMzkYvO6WpNRnlNcLTvvvEU
j4Bk5raClJwA8SenJD39avdQK1EDsWypfSVKqcoUKV4hvNOteWKZg8jjEi23TVRy
hjPvo3cKG7GDJVq3d2OOD+QvrGyW79tnzb7toT77hPe9uRwAxYuzFJADFDDSJ7OW
bpetfdbN5Dt6kdOz1G6ThxHRdyijRfGblA8NT35U/UfJ+/WfcFAOZ2IKPtgvmA9S
q0/Ozn8+I/jB1l1orE04LdVcgbJp5N7qRGHK2c5+TaURFAj+2fAODOqdAeFxkNyg
6KMQ9o1d8LadDJhH0B16EbVhyWgpTUcVE/KWCHgsc/+IhQbL6uZ5zYkg/zP31+7T
66jLgmdPUeE4GOZwwFxI6CsZFhOFNWm2ffxArnVWOiNhsJuhor75voWHUxba+9Sl
ouRGf+dQ6eE3/XE93tvPgPYZ8w6mbRZWC888GASh1hqdOERXVlZy4JUVLDcUiC0e
BEIKXyeRe+TCA5+UlN0nJwzkOHByEsTEXjJi1amYrSEe8PkL5Rm/eZ+3FcMqFXMb
PY/ssuUdH1iQpPb6nuVU0VuL2g6+QLLJos2yCXwPJm2jM/tCtMZRzsZ/h711PFEy
1B78JCcrgn/2g154FMRJjB5trI4TKRU8BI2wJmVPhwOmyh0eUrihhDojELfW25iw
vdi8jJDoDl7puNnko72lHUOzQNWiG914OvZgqcDUH6DxVNlJQllz6QmCLxyJvWCz
viCvEhguacIw/xEMivNIcalyhcgQJpiY72bfvJn9UEgFIKZJ6fRM7qhK9VXm40TB
tZtcN87kUjBxHjunZE8a4xdl19KMWFiVBGATKbew4ElL7FSTD7ufXWHSBu35EmJu
LtzvUGo6QXjBPcnZW3ZzeitdYah5Hij4xmUUKlTq4hdroTwPjyUHhx3v7CrkfBpS
6To4cwji+ZjG7je1HR9KsJ84Ep3fAtQYrL9epl+X4blAx+1CeaNDbbj+tfzCfCr3
ztbVQXcAz8get/M80skRE340Zp5CzNdcAxO05T/OCVdhbttYcOKOurVfy8JHRmxO
RCMgDBOX2m8i/ZBuyg4El+wcrK0nINWpz/COHejQz3Lmhv6HW/nEqTTmvR6aEMDS
ar+KMK2NQPZwnwxxYICMfzeIFm0pWmtyWmhvLAE46g6O8hgUfg1+qdB4jiY621co
0sPJe9gm64dnNYHltKSC7+c4/PRVQjqsS4AcUd2R24bu2iIsGrPFX6Rdg0MVkgXj
KWiBPD0oIjBAyT/j6DG09w2tEiFzY2pRzH448blp92bxuDorQauOWUjixdu+1zO8
2LiCu4lqxrO6wYkmMqn3lfTTphjAYm83d8OA+n7dm+vQNEHFSRA5SbkAeUJXmxjr
MasxMFWMpatfHaZnzdSXGn2sObRhP5KhwPN3FbY9qjafb9OuEIZaDaUE+gObPwbH
RdVjDcyzdAZL4KYVj1nNjfDh2BAiWkvnndQG/vyHGSz1z1Q766OLhiVoRhZuYbjF
4kv7XZy5GgdUGOa8R9Nb6u1OXO84XhxIyIs2wzObx2fTIR9fMYy8yriendld0eDL
qi84/bh9AIEL5OC26pH3MWugDYFwkqXaXIRJlh525Y0V5l0tR1qv2D2PF7pNfKUW
IUTeZgFWxgK4ya+ZFJsBNCYZS9J3AjJLcNwh9/SY7wOFeaOPXCebA9VXKhe14I+9
tPYj6/UBcnHaVPGa3Mp9SgcJZNkZDYPAhv9SzeTzci0lVLmcNwmgOVgY7tMBgdIm
DtTlfbaC6jI4y//6WHZhktk+3+lNbXBBccPEwILuhsoZb2nbPvtD8Xu0Ge0UlvYC
N8RUO7lNpDA9sQ12UK0fdgiQDEqoi5gGlgaiTWfjsRYv/NP1rzRQQSc6Rn2B184U
aPTPn3ix1pyGxKKFuT+ih4ilpBZXBV0z2aMUbGX4jy/xw7hxyg/wqwyoUjRx4EQE
dvQqjSJ84YSrxFF62pafV8PMmD7h2UJWcqAVCq91zJJTAvwSgeU52MmOjb+EPU30
VWzuIxAR9CAqVu/1r2/oqWPM5V05cdayoDPpoxM2WaECZoNbGyi7Oq/z/5x8Xawm
zLp48YFjojflb/ixbvvsdpT7LQVoZzRM5/OD6gatXY6xSJJ5un69sz24xcU/I47P
+as4sJCU+vEstM05NrORGQDQf90BCp7jTN+L/xPDcibYjfqLLk3ozGjnAVfP0L/L
h8OvIJTCQmtUnsoMGKJMnazb+0ftDa7fdsJRWDDUk7YiSNqqpEPwuYB8lq/lw93b
H5cU5rFe4TUKUrkqZSqoAjfa9D+TXAoms1CQuJfl8BTA8osd4wf2SGA9KqXLOoVM
iDeso460Ry+hT++le/7ZtqulOCAKCogGsiHp0Evm6SDdAH5SBOnBKlxXm2gs2ldU
LR1y98fy6eEqZscUs0ftGKNxOA+yJGjofj3SR/TbPGR9vi/vsawdf4llhiySgS+2
5gqlxZ+YM61QVrD4TIknebTZnXuHqjg7wJarN/t79jnDH7P03sbpYuHTeHRNFXJr
0z+TymWTWM3SuKueoZkZ6K34ucolD3bwvCa7myAjlhh0OSP45V1Bshj66TT3zy/t
IOOQrsGGR4QRbAVxHKkJD0eQDxmMMZyGUKcMw783PzWRoHCCrdlr1/X0av9aVIxI
Ovc05XQ3EFvSYVDwk+veO9Qqzj/4Y5YYjevdN7J8B6Qi4t8v8OuLr/i/mhz7pPci
0IJbxn4F23xiUjZWofGVtaIn7C1ACOUxyi7GVNzJXwDVuQCWK97GNxPPC3YfoO+I
HzQF5ANLQLLI8ujesWtgom71TUBqjUxScFbfVfbyAvnpXXLHkd/gqcC3fDV8md3Y
9lE2dYwYb1SIbOsaaxHgpRDuEvQN51NhnXvto0i28YUmaIgTT/QdBL16MOrdlVWG
/uE4XW8V9In7ZkWdSgd1WWvxIaYYgxXE6U3Qj7n5ehpGGLG/jUzTsawBsvLKdzeK
Xq0fFSJyDWKEuDZ5NYRkwV8wSxm26t3ZTybmy2VGON4SOmnBA/mIiZjyO1K0XI10
NmEsVDPGtsa0y1MoJZeYrNRs2DdY+xk8x3IDcZJ8X4n13Ip+HVlWQwOa00RIio23
V74KIlZrvS4znu8kkb4/o99u23SXZZbUPDbAUsTyZjECOVISsDI03KBPMC4Azups
uDkBozngfkzD9dBtjjhOI7VlZG6Xf7AC8mwX2EnRYq+rWw8mW59Ll8m4bw3tkJ2N
UkHdLuKskzKCDZMgMzX3X9yAykT1Kyz5bmsg67R2UEKozru96d+nYItqVoN0M6tJ
1oUnzWyMaSAPK9ZFBMXGlsNAVWM5bHV20cVYsKlBGnjOeMAcbhE47LgaZ7rqalFn
cusQCwcW9877QsVtQ+B7X3UupY2EdK2YkY93iF+XtCo/fXKpOQ1vIR5MuyMwu+QF
0BlM+N2WxRYj8woQbd3IZ7+Bz2SK/QAiNjch7JgQ2tQNPhx8PPfKiYJvMsbVeuBM
Nxuyr24lfn6JmXTyNERg/yZNQsm+u1sdg3sROr62p3rwDKH+8z0qvpNvMe3fR5Nn
Fgmsmoue4YuP9ikyMuGF6RVoWeF91+iLWaLQEoKPnnFj7jo3EeLTneIbP2MrUEPr
zKO4N9cJkcQCZAzTUk3rGC9oETCelj60+qDlju4DxBs0j0yXlVrrZSSw2tlcmc8o
fq+52OVSIsqny9V9RyJjpULI2KNPGuuSET7vpbbKwVLK0Mz9Z7fAhO8iRCE3KsId
Ju0JpFIJYUlymhsgHemHFNxVXINKQ9iUbHqGuuIv30giSXYHy08YABG10Aw2hrjm
/wvClMU67Em2xdsP+BXNrPZqunNVMjBNbT3ZciD92mCGVVK55t0GsLgQq81IWFSp
vxcfsgMYDOjH7HHD5765ZD4w475bdKkYhO66Y67clCBR4ZMs3KkFPvd7tKx4GGhG
jkbGXeVT5GnOUVVyHARa94LRuVypYghV6uxtSbqZ7hFzTMXN+0RP9Otrrradul4G
EVnKcS+8dUXbFqYVald2UFgZeoZ2PB6i9sV6JxGDZFpMSZvvWFH4+iPO/AShlvi3
BuOMAyDd/0KBSCfsrVK251bLDYMv8tStpnUY+ezuixBpr90nMg7gjrqqs4aQ3PVd
78och2mgS1DTKZLuoXSv0OWEi6rpKKhH4g8D1XSzKYCIKz3RV7mOnSV+Gq1jptL1
H2pd0bWJwnnvcrVK+dwndl3bEjeI5T/TN66czc51mW7fTeKBfzEl7c3CDqC9mTib
CUGaiTQgJLl8brwLsMXKgS8sIucYr7Nat8ec+BDUJTfyPEnmdKWB66hZcP7NLjGi
pg8oktiByR40USfBWlCe/4anyWPXXSdrqkC/HBw5fOJlMJxRH+9mYnx8ApQXnnce
Mi/wj2N+4PUWAiRp/3K/+EGS2VMs8y2EoLha/Cyv01XOGRfdwdDcRoHvEO5mtp0U
HiU+FqVklQV9O6r0PTuk+1UfXFrUi2QAAEhpxuXe4X6GSwcNeBI1r8AU3QZFJ7gv
vViSCDJ/dTn1rgljfRiEy3TUoUAPlTZKE4pvQKYweOCeW88NN3QZhP8iR99BDNYQ
plXbPQ9kXf0qPcHnPTu0K8tz4/opkVUfuTizkz1XWpKT+Qf/5A3ds+19W+MrTNNB
IopfzRB/PmlPSUGWZnucDQcJ7tRnlCCero4SYp633FDw+qrwPQxxRCCbstVFJVLv
jrnI0dxWKg4fLgsiNdI065EZkwL94Ov2jK3zasfJpDq+WhWyHNZToT2sTOG5rIXm
7GsPc7THuBm4qWNN8lmZmkBzYBlYRPykx38MUTU3/YNcwP1M3dSuDpgLwnrk47VJ
7fP9Q6xixhFSKV7rFb0re6sh5bvwN6Py8SYBlOOu5kG9Qhx9wc06/An3vXh836cd
56ibeOjpPC/sYYCTXYDQz9/cQ5weFAb9qAu1GImMK+IyHNH/7DpoqcYP6aZnIuKa
TQNByPvj1qyOLVbdhteK3MVyMQJzs9xBQDu6JydXk6fhFzSHcUA9Xl7YGHLDjB5K
AVhOHbiwlPvnjIEvErtvEXaVxUxnrflea5K0e1CzW6xi0dl0YbHsGstk8X/2Vz0f
QlnSisY22QUuu/M2pqrM8MPtnSC9EIZDbY/l6RqozNhKjfhhZ2S5xTuFVdiP1AfN
vynLVbDGDylaL7dTlA/925JnAuEYInXeqzlBq/Ele885f5cE5g2iji7/3uElvAj5
DJ2AUT3R58SbaZ0dMLfcY+m+ZSVz292UtPz1rKJlpl7GoO7PdsoNr+63P+QheVNN
V8IiHwQM9CErpQwdGl2BstbMaGJzoAb3ylxRDUWLBeDPj5Yi3j582JHpI0OVSOs1
J3SjnMqilEJBaFY9jkNFTl9RWQFDJMnOQycF6K7SU3qUJ0rW54+4o33nwWZnjPXu
rc2uvUC9OQxhmG1j2ZjqKfxX/A3IN9GnmouNWX8PiyaTWXfPR7TPdJ+9q+KTMf8I
d6Q0zjKeqadOAEQtJeWkY3NwCX19Ll/yikLPE/LuwmhCsTwbqQuURsOFl/KvWphY
J8ldVvH1b3BUAHV2ndpwGP74G+vh9eOf0zKAalucR/DT1FWU4+IgraFNxKmwG2uq
rfc13M0tJ6mnp01HXzfv1daWsKHmZo4Xq6JnoEWAefiMa9/m2dJfdDc5K4ri69vu
vAbnl193mTPi7+ZuTp2A5smuufafuoDVWAmbI8SGl7nGnObdokYH+rawzYwRvy9v
hxNx+NiW4yheKzhj6dH/nOUe8cUsDG1+QCM9AzhWTkTkmDaakC13bSbqQOyAsCl+
e7pCbC929zdCV51c6M0n+8D4FJ/bZu5cHY3w4xbC3UToO/ACuuqBY2rNJqFp/3tT
EacDxKL/Iw4jpLb/cweQq4PbWpXSyeZG+k0zFaKLY7wpDnvLaLmI3W11qKaMzRE/
torbMcE2+zshlHDdXKTw+ouSuEA6xRiLGbz0Tky242qLMcD9Iq8DQKQcoZ/puMRS
ZrlMin+ue2Fcg84vLGzaZdU35AOd0vg9+6BJaCRskhoUqmfCkfCOkrVZ0TSwZ6Cr
u/Xobl3nmrLToQGHq5X6s95Sh0q3+dUoF+33Z76f/fHwRT8HDP4HdazJbHd7J+Y2
ChCir0PS/D3wrDA6w2lgAxX+FG1Te0pcxCxzGUMFEkE=
`pragma protect end_protected
