// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:32 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CGzsznvctZ+2syiNmxNh47jwzAf99qn6RkeZ+qQNAL5DuMrNxk/Bw2KXSRUF3lP4
DDCXkSYM3JwnzNl/CxIpd41z/QFbgZIdSZnljsOs4DUHpAHnnD5wehD+yD61xrr3
Ksf849EFLjN+1aZIEVTl8CtNEHCmS5PMr7GNohlUoWw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10960)
Mcls/5x5clUsRel6XvKDSFgjo6aZkPLaC9qvhqTZvhbJHDhw0ts3rE+Zw7mNOmFG
Rc8bcRoauT+R7r2QfC5EOQ8qybPTIbGtgpPw9ncVptKImtpBfmSYm0VQyQ4Mjg5a
5Yd0Ju4hAiBYvBL9qUlXN2wtmRowxo6+7iazA0zZh/+/hrbo/fOZkNcFi6m/hmj3
LOZtEp1wFJ3PpA37CsjWBIMmnGMBeCHcjL8liOU2uzuwKWORmn+eqe1f5p5F6BGR
hbpzozthl4BsGr+tup0KFBUsXik2HGoGCjId3dspji+gtST1qUUGYD1scbX2xyEH
4OX3lXmg5ETiNmZ5+hrp5380yU9+NNUJh4EhZBi7Qn/JiBAf2/CUqA88bk/aS493
Tcxmf3C93TCLaJDB6PveCsCHfigmt9bvwxXn1iBdrr+qca/jQ1LmoaiiTCenLzB2
gJ5QaapBY/gCH6JtiVhnXPvySwU7sYt6xSCo2U95zlD5ntLiexmbQr8iSesw/3PT
OqhkkUExZJ3/bbap48yueTAm63OUn6ZHyakTs9FlSLstqIcoPHk3Pi56iQCAL8tz
U9UGhycoev1J7dMAiMxaLEaQWUECxwYh08cPEPl7Qf0VGpMxM5gyePOhoBIm52ze
BEDw8hs/Nd3fwp9544Itt+6ctX01ByC/70sIzcvWLmR7C7nciIFiVsLctY8D4LKo
vA5CQDdRLTB1Nra+tuXWxlLnBliOxNhpOvWrvkFr70ec5+/POhFshbceG/fUh+Ct
6nSCQK6OUlzsCbCzq2uc8/78Ci+gfX4i/2k1/UfeBoy4vt1PlFkjnVF2EHxDdR0P
wU4z0clo28NG6ihuRXqKm4O/n/HMyHEamXGuJ6gfD1XhY4Nf03NIMBD11P0bNfkA
3PLkA1oi/Z3iGJ16I6jOVRPCwm3x5JkeBvPyLlJuNARXwwkbSq5HgMXpy+fmEfF+
1sFMdp+aWTUPkuArDuZcDokGgNrSso102EU/ia/of6TQZType6DCgxsG8mTecV4X
slpAawZtEnayU6VDLZR9aroUif+lSnz2dihJDufSBLXD+Q9DYQzNa9GAbBdXSjAb
hJqSpvxafue9ilmnsJU5lDlXD8MrlEVMaWUpdGVbpBj/f1r2IWW4bfeSMXt/XhQP
gfuxyi6u3CQWpAEsknGvrwsWSNK8hfo1oMv9Hs9MaFyv+SiuBJmb3xpQyOH4sXjI
7jfkOdXoa6DQs2eLz9lztc/Eu3Jja8Juqy9ISO6u8c6xanklqDv43G1jVR448vtf
Ta+w9NbxEFsMCV2OIb3pYw48+kEZzao8jOgVwuSendylhaglo78T99Jr4IN2qadI
FpihX0vdoeuE+Lc3UfLYB1rzdecGyS/dsEJlbabzKR+yLqn/2mBLwrsGmjHjCxlM
BF/VRP/OajBJGYRS4/tu7rHGyA+/YXNIN5la6Q8hKIu1vN0YfP4ag4i/LVZ8oC4U
iuVJ2Mn+zn8/eY65A87KEXyd+gyH4SD9R6LHuzJqfhBeco9GPxxOxcs15XaGpKFe
r4CJDbjo1dvmAAyiRAZEDp9pvtY8Z/QxWPAeaahv+7BPlD3zSgvL5JCPm0xig8uJ
+8+iLZ4Pf2SRYD2O/GQecVdFsCRgg4tjvEN2w18Dg8LQtvYonmuEWU2mKUYyPcde
o3wh9bW/mOXXFdeCtxS+t1mijavr12AmoZ6JCfXH7ubJCUgpt8igA1MXauPthcp9
PcgV4wQbXd+FSzJ/ku1Rj3lPUVu8/+P63FeJzjzHAywk++9aeDemEttYi+5nNL3/
2bFxWadhcGjF6Js+3+DYqxEriHfOExgC5+DI5f8kMmds2s/rck0MpKqBR0EV9dOT
uMRgESrt40edlAGNgwI4qKIjm4T4rwNUByg2ZGtnYwZbHR/CtEciX5rtJ5poTMVA
tJK94G/lTkL3zEjTA5sbf34l7lJ68QVhhFbbrNx+7T2VOWMR3dmmizHAgunLuhMe
CgqrGi/FplWAUjLgOYyWN3kWIdIhJD0+VXa5wdONxYh3kvCeOrFW4+rTB5Rolzal
sJXRdMJQBeZgdOwclAl/xFa2SW2qC9A7EOq7NJJwnvLiETvgKwsZIVvsYTU0Or52
I2JAVTVhMMjtKYSTB18a/AwOeKCiblki1pBuL5r4uxrtE8v4i9o6H/Vx7xFksTcv
evL/xuZN9IKMqumQN0+DHSdGZENtFribUyeb6fvDUyMFdQFhqhAJdsR7NXXJh7hY
5cJ6tkLrjsBwTaLAEbCeg1wYUgwqmggK49uV0NVicjFXnbcGoguo4wkEwSCkVtYy
TE78BjTWFFs0h9XvuUOyUq8UfPqvSAF19qVrmpSkN7JPr0oubGGN4ozHnBt5tkj9
ArFo17TCxa0ad6oVAcQF5JAngSPxhcDjC6m7rVG0/0QKhqHoe7kJ3YW1yxYYHsOT
E9JfTvgyHKw69LPZLerF+hZ7liA6dwoDWoiLZL4idQ4F0Nspezhi5Lx4SunzqXub
5HtwtKMd8eSQiqTYgLRUZin5kdm2/hRYwFNgUE6JAV7/CMZouRp6Ke6dHNFHQvO4
ytIssNYAr+bHIxasTp3TRIVYLhzeFpcfQ/4wD3uoxotwa+nB7dNOFxPMfh4N+qLL
CDMWoDttWHlqD9Roq41TTIP149PrtA7J7z8kfQw0pEiZnOlO6FEX0rM0GdV4qgiQ
XiXBkVmmDnu9yV3Kh4nH6hRmApTsdD5Nb/UKk/00ZV6ADY5lNR2kTXJEoz9y9DYr
IaFD9gHJrvliypyjnt9DiSk0pDSHOoyyLwGrHj9oI5ea4Qn17Mz3SeraY1yxN8j3
lSYLGeKRJQ8sgQaJbEpF+gC+0QQI1ZsUFf2a0ozMsw5iJ2xr4OAA+//eGPsyi2Xd
We7xliVEXcX2wnYg0kywWpLPlTII8yMIB6K2yvfC5dOMBDMdrCiZaNYYmpCc5H4H
ZCWcDWOLTSqTvlm+v3Frw0gwFqrq8BY4/BACw6OV85bpmBAcCn+DQWCp5UMjgqOu
7aI3IkTIOgbjmiq5NKDXrJ8Tu8tAgU0H2K+q/W/rzn7FM7rqsDnbNAL3RVnVNgOJ
mke1TmwAxAZF5UJ+ukhROch3LUl6uLVbdG+/Oss0hfZMCIx7letdK/QN8wp3kCek
wZYq/Q43krGoujDzzour0rTbHxhdB1tdLrWiCCAEuXPp6Ulz2J2VMnxK5jk0Q7or
tc2oDror619k9srYLcmNjds1VorRXjW1JQeLsjMlr351ITr+07sd4QSyqJ/7P79r
WbCXJ+8kpdfHA0HlQqXousY19DznYraEsFVCshf+IltLtBuCxGkZakqjT7HM29fZ
QQQZaxAwvTKJqqoaHLJzU9j5QL+9bq0ez2H3ayS/r7XofCbiKDsUiiVxgsjNfxr3
fEHbuEHAj1P6Pgzl3+ffiG9iFZDuyNs+FMGFMEC2SZOyiYEl6g8dYQXYYbsmytvw
T3wXoeGfV9TmageYHILhbF05/zjpbpLXZaylzBjwZqsiOvTeC2fMgfp0wBBnEPiH
QTqJ6eKr1jtdO9IOGTAE9nub630mqRFl3BWr4Uei1C6qqCv70QcpRsjWu448D/XL
aYYhYMWpN8s9orH9K5LEZkgM+fnY4JYkFdhnwxq0Mp3Ypr5raqUMwFFBJBgpZqsa
DIcjQv0vCEG5Cmu3xqeChXsI+TmiwiSp7/du5VEfM2R6zM3Qste0qHL7npq8snfL
H95hu7gqg4BjkkufEUDXFU+Q1DCJKdCprD7vCSS3jbVKUKgvHMhE40DybdQxKCyG
O3n8I/22GpFANv6mSY3MzVq14lw/0chjsBKpaWXJh1ts7I8XWZmMSROyoqtXsGzS
6cWgB9Y8FFghF4YOxHs0D3bjOK6Wv4sxbifTYK3mxYgAQrXXjlDeZamgcP5XKgVf
uUAZkXfNyXtweXDSsW9X1v5bDt0VP9DKRBHRY8w7SJ8HCZvUWGueqDhj0M3CEQuj
i0Km6bthvZdXN0K3e7HJRD6VlIpNiJ8h+Yi7KJfKOEC3O+1Fhi0+uVZtSVn8y5wC
j1BNZ8iUulCUiyOWarnWQySjSIyCNvIvi1tbcWIUTuQYcN0v7jHZLIt63Xt7y6Ls
1ZseAe1szhmsKRLa7ij4S0LJZFwAiCgz/0LKrbQt5lcQTkcp1ON5xN+uxeqhX3vm
m3wcEIRIdLO2yRlKkwJ5rRf9ED8uKf90lvRjFs6dy40457M/bljIr9UMy9eaZyNa
dH3N0yV/8bTYYJXLkvGRNTZWk9mrkBujdRgX3dWhNmuZ8o0E2kG+i7J4sKgYVjig
yDmKzrlcKzoLefiGpB94h7cYVkvGhixB0KQUBZPM74o2QKOOGDi/kOerDEJlcv0S
2TGJsdbvQvZMHoTUvBWSu8iwMzM8xUOha/y7P9Dedow/2oTryn/Ap+uAE0Lcu3MW
5yguamaQo5UkPH7sJMZ5fVmElX7sjnMo5cvfXnMpDxnVBBXuU4BzLcJVUW2cqFDm
079VgVqK2FlC0X8bfD8TJ0AM/LK5khrEzQ46LUzXcwcsQKmU/mVlrCPFOnL3aMgt
DeLQjm/RJPo/MkJHtSC+PrdEg8qJjkwnutBuieKzWa6BO4mWNim0W7uGMI8ckBam
xe9JwlH6mGxNLrF2/58ZlNYJvSQ6PbtHxN5ZuvIX2Vu+am8eDXxGCXeI3X98kwdF
qF4B/mlooCWH4uraHEls9AsX0m5VCXxXC2z9JjViPpJGOWnB8cv7fqcgqyNmIb0E
Ig3vCI10m7avbE28fPNqmUqqXqJ3hFjeL1e9B/i40Jc3VBiI1Z/GaxYkQGIlHRbU
w3hmG0YAxVEjF25u/ckf6Phf5zIPIOSFMBnrzyOJzb7ZT3+5aROYbzeB2KKrGGhu
N0irNdmAgrQzsFGLfsiiE5PdxeX6iePtyTtOqYgJJXJ4/Yj+ugn6IhIG+BmfqTJF
qFl6Cs+ump5B5rhmRWxLwieGUt79nFO2LLjkaP75cX4WKa25nE2v6PvRTNR64hY+
/g7kG6/w4XB06UBBMjgj+1IVy3r4tx3P5ZGtWEFvi4MgT9+6twO2RMMcPJPwOnhW
WvQPTSO0XHSoe8/N9e52L5bgKFegWevziLE63ybQBd9Z1cwrid9yMjKILJHWJRfM
G1eAuGnmUkpKD8Gb8kA5oJCwbNy3KkC8zQ2pQ7JRwA925raK0/EpVfvHbULr4g5Q
5rAdqlvAfiA6TZwFiEEm5VWGj0hvJvCyN7QBikt9e3Hakmo8xe68UiRGZaY6mMFj
a2D68iAT5c3GNZl/yg5QdRujn030dT69JAQmUXokkqTslETL/u1+Fgtw1Ugp+BDE
7Us+0OZwGXVWq7QuwHFDCRRK8ky1sNT87VXRSqBh6rlJCeDyNrDIwolOCTdkROme
OBeWsIOoS1VxgXn0yz8A5YkpvCP22ekP9QM6peyLrd+5UMgrHNJBrLu02LkNveaX
7xVpeGOnn+1vPvc7YhKg5PpVr6BdTMMWvv98OBYNRo9r00lgJAXINHAgfXPCb3UG
3vqU9MASL3RG2Ii8V6Q3JGuhe3WrLnp7a++cOScQBcjLLZO8Ui1RblGZSZVAFKXY
ZvUsd7vLfDd+I4RV7ZUCs6AF3xEshioIKKcHcNhOw5vmjrELnNCdc2loJ1MFQQnL
AAndT2MS7VqN8EwFfUqqo8e0D0LwP5FjLbIk0rbJBrw/SEw7BA0NB37Wob637keu
mjCxTY8b00tZN7uk3tPMCye+KSQF5oTeWYj6XyZI0Vm8QIFZxw6KX0d4HPh1R8Cp
fc40fibl1o98PGvCbBxg3qDj5T9DbWbHwZncVFqtImtMDlDtTyWK9x7t5PowFVoE
IG22k6HqESTC9WTFPj9J3QAAqgJpuOmaGV6id5i4JdjOBdwQ4QM9gCHa64LqcDtc
xrAMezpZTBN6mxYZOkLjX0p5WTccczkM4V2+jkkSJIDarHxpdrCzrhtWGzWcBbwa
LZ5qeySlQkZiP44VGsxtmMw1qde4K/CJDl1qyvjfyEnRjnHrd62wY/WNIvejBWVB
rozWNacQSY9BaxdgvGFzM8II1LTFqrTxssKPAbXWSgfyPYbp+4Pf1FdOP7pjQGa1
8YmU7YMFientEOHQ9tNl38o9yMtkFlja+58LXRYC6LCm3ukf7MmRGCD2NM3AWHXa
CTGq94ByGLSlbTuZM2cXXUsgBOdzIPy2KLVSW/DLrrtcpDUvBlzBLnSOX7mzApuV
iJehDHYNKe3L2d9vIlEB9XOSF/XKB57F+aCgX7hZ0t0qDYuzYIQmvA/JQNt/nSzu
+spQLsRTARd84pUMLlT2tXndFvhuEX68e+auLTX/4D4mR04OmxlhJSlnkVvZE2se
3iM3AaaCPSddukoAW2bsixrnWHmHYgxnE6JlYtb6/SLPLEf+KfkBLYXZCYxXW/HF
U2cPiIEal/SnjbpKu711fr3B1VMBrHp7QIhYjXik/umNLMhKG1AhE5j3fvjGfP5Q
1gPgvO2rOoTm7bhaoX/oSD8sDjhyQW+URtuWpUBPXJEw2buZw4wuJ5XUzhwsVEMl
omG9rGMFgJUtohFx9Mn/VXVwdhbRhvLQK6pajEdlvp7VSyLqmwcvJWa7jkR6+pJH
sM0dD98H6tDwWUlliBofNQg7pNbxrv9VQ2uKCC9JIU0/cAE5CrMcYlrivec/LfnF
QhOhh+jhLsQ1D36ObmOHAM86DRKlF97v5vaFS0sFYilYqihQ9K5voyPDZqIMN8/9
wiAVHF6r06NU2eaqiqCSgsCy4RDcQeWVi07U4VRVzJ+w3VG+JZsoiLgOqWWVCIE8
EZI7xWPpwPEpTayFPMVG/19G+rI6plAv+j2ur5YHfReMgkch3950o7y8g3gCkiO8
fffABnzBfXdUMf7gkMhdsuivF5eqcBhRS25B27vejvtJ6wmUUEcbKJ3JjybIgJci
v2ceeEBlFiTqnh1wjambfUan2kuc4sDCHMGaBmNEPWbbv34T/1h4l1PHAYQCEVgw
liTZoht0OPaTJDhhlZvureLVTbanoMo4EtS1UajwZX3l6TS7GpLczBWnZ7m1CAFD
ebXqrxc6VSIoM8jdaz/9fC7ZFwsrjcGRhFhWQgjREng2vyMjKnM6XvNgn4JsrBk9
DXIl3yND8KpIL0248baHY4W1rZWsSIldTGLh/6h7FMJRWebWudW5wQ5aCVYllpn7
L8XK3tWeEQnk8mSyJ8iHlSGsW9CqkMvG1OZ0/DWENFgNwU4l0jpuNcv1a+UGQC/y
bAktxDgl8+kk+rQecrM1q1s7f7YWQOxnRU1J9RlMDC994Cq4uF5K8PgB/sYBkFIs
8QAb+pJo85rZ4C/p2byf9MbMW1P1C6M9YwDuamFVfMDnQ0r0FmI8EZ5ShctRHCdm
57Vb+LfukTxqAR92WYFUSYPTUtScptjYdKSZVyILpZiZgQqAHgfuafzmRGBNXi8j
PhWAoiTeuysovALEalLzy2ynRrDT1js3ZQMDxJEJC25GvdVZLCtGjc7JFMHWqFuC
aDZQEQL/sDLLmSCgITU1SffkUwt9qOHuyRk6jcncXylXFxfhzTeL0ZxvENGBUp2P
Nd3/iXGofU1Y3kOg5gcVUP6cluilXpqjlW0RYQ3rkNCLnWpa9MttflP1mrTWkJHV
QkUb2QW3AWEeFtbtbvIIXzF4xeu7asdAkC0Xq00YvZb+TUxgdgavPJ8ITBaiISKC
x029/L91s+B6RyvdakWXY9zSjzy6klk6VTlDAUy/vfCozCQQMpz6mOHRFQTEr+7D
y2q9/2lb8DzpBiTmx7SwElnAwOiOHfiPk1ryx8bkGq8P4G2ZfxCNnVsA7dPEJRcO
JSjsmZnjD4jl4lRnzFkeNCkgJABSYbtxcEBPYvZB1J3Ik9w85NWYOsTfwrR2ekoG
xXoZHHej32NWf88/5hgCbI5ooUr0tkHaDET1VkPdomaczzNTEyID4Z4WbKp0C/pk
kjFpBGAX/P+e+WxJH3+2dgWjgHNdQyHBhnejRecfdIOXERudCCk8gYzHhZPI+BfL
YkEwfPagiNO1cPiFS3N//0MdWJ8+Supz+OYEueyMH19dCmJ9+pcsv8x+Imw4Y1Be
3OpRnBPpm8mdD7xhGQZBlnGz3XTaHbGXl0IfuUsG2doxU7Fv6KmAt3F4iaONw9Js
w02pGGtzNOqTTBbD+4QMK6uEWFOfGEUAgDP0LZaUsdvzZmwvKU71nXVigTVURjX9
nE9LiCuNcuW8fCkCfq8MMAiS6/7Wvzf+82VuMeJFwqdFbL8TCModq3LoaRbeFIro
jiqcUJ64ukeAMn9zeT2yRtn90128IMl1d0pl2OMuWn4BEq23YFgNBHliw5UeyrFZ
LjCsG/rb5jRGb9nzmULEznXCmVUq6OzqhHsPHh+QRIHavlpUvh++4+7Paf4NZkw9
5U6v+oBLAn4WvhX957D4EiYl20uRXnMUBMwAciV2n1/52wX0HD8pURoq66ZZNOlu
IeABL0yptLFy7FqkaxCqeAHHJJsf7psNYFWrdYX/Vyo7ZHqg7uB9eB5lAqELN9xv
xGj3jbgJEGsv8qqzXX/zbKs81V02p/0ZNfebHQ8aqghuho0wCT0In9n31+AOIrfK
JsnUQ0Lh+4AZMWIW7TrqoGH7Mh1O2NeVi56f4PEwZ/ezCijJ6oKiZX5lQ0vLEwG+
0H4/KC7T4Ie8T5hfaVHMZXWc6HgrAozCSSsdib8yYg9P3BHAsno7foUYiSB7yUKx
7pki+LxaeHJglR7cocUFLLiNYNjjMgQrbD7aXaCfuOgXNIFeUEdUd7I3lmL12fG7
kALkUdCY5ajYBoea5fngMwmHI4VMhT7/jQ8OSmuhGLUA3j3N+5o5aAXW89u57rFV
cPeCRxTHAPPvu+cWXBFu4HroG4OTYlxPOz3ml0JjO3ZJ09/syzpd8ZELIU/VOcQZ
UB9YZSdxUi4j7kIEjCc8QmWFkU4YPho9xBnL6AfSROi0QeK7AO+qaiKSTwlmZv7I
Ev9Pu0UT9Pf9qBuXAlPQgAkdJzzdN78lR4Q2ZKvSQCSos0uEkBoEHHgFBSGTTSE4
6bN4xb4EfMnHVd0VyHssce34nPjOrFCoz6GxT49Q2TbEh5m4DAS4hQX75HWAPuZA
FR19mUfcy7bNdpWKjKhJrTPz45h1hyFdCvVtdqmFTPm+6/aNRIy6fC3FNHew80jC
pcj7LwT10OZ0Rk55zsWPZMJE499lHRJSAyKNeWDWvMEBBS3GfQZPFrs8pjBF+bBL
CKaJGbNRZVCxCb9mp4ZwRe4lVomI01avKFxJwyHzEaPS0VE4bMC2p3KGZKiuGrtv
r3mL4qMwsbRZPPZLvJEgchBOviyv6eblvXi62Fi1auUUav1i+eUM64ONNE26A/w7
AB18Z4chspzKSVFCa6WBsirL9aEc+EcpSaZgMyPipsiIyvvdADB8FZraW1ynPUv6
n81P5TpE5G1AjivHbzgfxTjn8YzyxT33/y0r7FvyAE9l+oS7XllVVud5fkHWYZeV
cbrAWDfAYE0fOX2SY+YvykC5P80Zuj3Nx2l6hunJeXUOc/EZi+FdccpjFyxaButQ
yn42/Cif2e5VZqR1lwn95d5VAC8ou8ESdDgWv7qzjc2U90kaVXLuEwIAFHIWQTGK
sbJrYP3ByVBkQPjQhOFHn1vcMUVU3GSveyUpv2v1yiMneKB9nRPHxbguUnOUWiXb
1AYPCx3wzmUNzuk0i/iCB/X32z4DQ8C4/ROBL8sy+YVnRtawrWpIK0kz8tyXATc9
raIao5x7bZPbismxPcLbSkVTSHltVTDZDiWp85z+6+FlKVO592xa/aRJjLL1tkwv
tmYm+ip8ulIBFwy4ihpvqiTTbVVnWUPUQ97askYFO69zQlvNyFnPE33qvBqDszJE
p0ymtwoACWUd2LSdG6aGRcda/dkvokFkQs/Q6eT8Fa9xzK/tFfD2jCYAjiFBc87a
jdfXqUDag7x+Wn9t1SQzvuWWfEodOlR7G13INVs3OM5A5duFTRPwa4zHUOut0vPA
2nZ3o1a0oGzNM1RPgoCqqyNn9+gxrVl7I7d8xstTNADO7/++yT4x7FoUF+GOHg/m
mOAEXlrRbMgazRpbDjuTUyY99IH54GD8keL+xONx8rusAP+FEgHRStHxAxZj9KhM
lbGoLoyogTUWBqq37EAX+Oh7dTBEqFawVmj/e7DIEh3xNM9sTT5upcFlV8AEpkPr
/CvthKKdmiIfI5zncGJaSOfIFAjh6OAN6ijqv/FM5mSeTfNPOzbt/ZWEEsQuJbl1
Iv8hLjDyUWVIBcw3//5z9VE0kmC0TMU8Ee9fr25OtrcQnZ5Z132pFu9BpFZCloBV
iHoaY88LExU80CqWNydLNC3v0Kdx6mgZchhZEdfspc7V+TMR81rxXxl5JL75ahig
4rPs9Hp0C7l07TQTf0He9sHzO0YCkelmDZ+lYKMPppD5lbsQwme8tHKDnyWBud2j
DxWtkE1+nu4zfHcalsafNB3BEN4ssuDTWlcdOvXf+Y9LRYU2cOomoZ5exldl3clo
qdpOp+MpV8sQU1ocN083QYYuKHr+prsERj5ksDg6TYeefo7ShEUjQ+A8XmSRAnVT
LmPMyHVY2IN+S0KuaG70yL7YCH02r0VYUk9eXuZACIxkDKlActc1jdrM16h3uKnl
GcLxVwvBbqlCY5VIqgQBe9N3Fq7e2mGRbMJD+mWljomBeklIcdKdNCfIZLxAxAz7
zxd0JD7JmeLVDBI+BuUZE/+TCNUUnOUpVV6zRO03roj5/+M7n7c1iIh8/fgsNvss
E582A5qxZPEUfPt3cI1iooVX5nB/SRDyHxsXeCOdelkTXFGLxTYjks230MVjydsd
hEYwIuNxkD7wExXco4F2dVXnvLSbvfDwaVIY/DU/fBYIH9kyZn6YNJ4Ql7DT+/xm
2LN6HZPZbTxlkK8LSO/cIEsowukje5CHFtZF5h+rDOBFI/wuuT3QRBr2lg3vuNjJ
dDlcCf7lhWU+oZxiEBN7Qo1FM1yGEFQ0PgPznwBWHfgLzb9Up3pnM100ITi/5hW9
jF/UzYG2bY6BvBCqp8FmE1opJ/pXQh0/D2glqb/YJ/ImaBT+3qKb86jHPy7YJpm1
tX3zSgqhoVEZMX/8k8x8gx82Axh2v0APcdYxHu6QqUEvCYhsts3Cp8so3/0HZFxQ
d3SCyuZfAJV4gN0V2GN8tOEiNRo1/KlD1ZFLd/MXKqbnLQlTxRz1Zv2ImfQ+CKPE
OUYx62PTYt+WFldnONlKVqfRMR2PLudToELgYV0Em5/rJhfshcf6PcjMrTkU70j4
DZt4cj90v+moGpOwXwUzwQi9u9JgprqvT/1T1MvohX8FqxMa+g/2EBApQwUxlTSn
HP1oCB9K7XZvyYj2WyzJUOpMoqomrVvX7AF+mZAE4SVIm+HNKGZt036WmPTc1fgD
8GBqa5U8ana+AqHwB+7btOuviRy0xg/B12gl7FUvSNHM8i5ETABmwcu8d50sa6WZ
Dqqk6S6USqAQebzk267E1wmftM5B/2LslQH4fSPC1sIcIBIAg4M0/rjejNVbGQD0
93g9UIBrdBfmMU5SqtAchp3vgSBOTOxJpT6lxBdXklbeknTxXAImPUvJqaLvI5g9
UAGA9YeVCuUB5MJYUIAnkK+n98zCztyxDvGfprmunMFS59nSURDHV8DxLDidliuh
yATeBJrR5YEvFlPti0aQcn7ENI0OSdD2FeO5UJ3u1Sa1ZDQ+StuxRMaAwhEwB0XH
6wkbJetX0kqqz2wg6stHx1f7iltgItMtgLMMnOgMl5eA6+Cgfm+6Ecv4VQUN1asL
WQ71dXiPlZcsUjV5J4sPNbt7u78+frrP9PysJ1AmoocRC22b6rYUNZ1AE+WOhyqH
g/uVVFOXOfaVWOdxg7oeN4HnEYUm5jwRY36FBfG2hRY9VHFGPJ0Ov0IqsCVa8Cjz
KdmSmKZoA+/PP7OLsD7FTTIauvr8tVKm23w8+a01/uPc5XXEAzgvM5unOkXwsKrb
mXfAfhvcV7TtxIw1p8ujoyXeqFQV9HukZADsQHmOT9sfpP4LCoGN4miEdcjPIrsY
RKqIhBWUym0yjG42zefBM5ZJBdDZkFbVbjqbg2AndfOUdDiV2llxPz8Pt3bPwiVV
GYIsrsEmmVQpQjetCBPxhqUpexqCqgk2RLu1O3J2epaYvSHG3F6Nv3NCXw1kiy3S
kxsdxsdb9BN/9wFbvQFOG09YD/euXdZm0qQ58gNYsf87FwdsB2UG7hMlSH0YDiNg
eHZ3d13WHrtuwdfoAkwBHkfUGL7zd/KL5LBoMPTb3oI/xioNHus+fv4cr5iUkBYP
emU9xtanUf/JBjbyfo2/HgxozhUzVsP8HXOdgZWxDu1Q0M4qhar4PJc38oofsKkd
tt//37PNIeEvuBzQcE52N8sif7t0AbR+PrtfFs0JBhXzTmkGqeuBjE7zHa+MdWEu
8SUBCaLnYIHOgug4A82kzgpFMNtGSYo/GNh8WaKhiLo38PcnvPXNZEn9yraQQJTN
IkoAQuAmpjmF0Dl1wO/PZl80+O3odLIdN8ugIPZzXtyAS6iqs8SwC3lkCYzlljIO
Se2tmwjZtqGVdF4VCn2UOm+ChPoD0TwrjVLoq1DwIBRMupevUb+d6pN5x/4p8d5o
YgXyH1WqyLCf9sZYEvpYsEjp1j1Hvy8BFnHuujFJ+bGzo3MoHWzIZzONaEkj2i9p
8cujYykt928SdQ7VCCeVi12AJzBB9iwdRV8ivlCG0muS7W/riLhStQQJ1JhOpQVV
McA6PsYX93FctvGk/CIv1yR+b6wC1+oGN556PvGwe+skafzpAmk/t8vKLv5w/FyT
FdGguCihWJYN1d/CwAiSdhrWP1Xnffo2VVmbcpAvMkThdwa34pufRkChe3BrNqu4
ithDOIK0FKVR0LBcv7w/7f8vhyKH40H9hBqYDxZY9MWho0c4KhN3wrVXkkd2IPmc
6FNp7UdZRj0HcrmPvNr69oYWBM/G/8auT5tD9NmNEdMBU6B+GwSUGv6FWZcU/W9Y
ly5m8duyF4kkcxTj2LCaidFMnC4/Z2yLT52tLpHwcwAWngmD4BqOunbMsLJDiYHg
UJEuL6Hay4R3dsCYmp7V+65TqMqxnEgV8DhZveTOIp/pt/YsGn5r69/YZW9HJAsJ
xLu1P6w2t78iRmBdAjm2eQE9Q58yrThzCqZv2B8DZRid1RJzkDzCOq9/rbN3y1qI
umdOvHp984DezKsWdNWhSI3sN35Z0AJ4yX5Zm+EbxGTi+EkLI610kpYfFqBKK93P
kmV1elGNyeBicgLJx+N+w9ww8VjEAHS5ico18Xv8hIEdTUhWoHl9IREi+f9Cpvuh
kY/DRvSiNRAj0cRo7W/iTPz/LgPFRx/VT4oOZo0qsVVosAClHleWx6nug77lxUB7
g+XPacD0LlEhAbsL4bISq5UbYynrTaGaLkry3u/jeQ6/tX3tCVjZJIhaX8Imozfo
zsWJpa2b+DtMcghbGEjCU9o+b6U/hkQWXT+LySjV12GqWlcvw8IAJfjOv7GOLQkc
UtfF5wc3gfsEDxrUJHSFNPfGYVUabxNLJbn+pvAapmT9VjEUTPzk3n/R4VzsZihg
bpoRGt+LxSeYK1YHImU3kcVhcLOG2n44MaBpo9vGY+upNwELshgyBnOxkXvCW/M3
XthlK+O1fPBI324dAEQGwSJLALgpgyZqHwRdoKyO70WyOE5eaYTSqV1UB8cH16cX
4kdiuDqbSGTF4RXpJ3vxwSqt3om9HLZdd/27YljDFqdP0iKDp6SzlMMAuEMAjs13
SfvGt0rPAm7sLQ9cebrl6Ie86MkezdbEn/qhpo2FtjXT6Yil7rCkfb72oryHAd+0
y213cJ1iY4cw5LFzbX/gtYlUHIk1sDTkrPWUNDv1a3cZIpud8iE0BYz8gbM34qwJ
NhhN/lcrzg8Mv9DPazcKtM5NR5vzpFa1Hjxa10p1ufHu2pyfTQRDK9pFpYjLY7Px
5Jl4GXUDt8yOmS/x6U3S/KloC2dq/CWpZs/i6lcQcZVNK+eO3Pbo0e9AzTBLKdb1
QPgsagviv0DIAQjhiCfLkex2jbiKxcAncaRpFbqv0Oo+W+NcdCRAuaRX2TRhlmem
/fBq6VH8JesM3f+KiZd6OorblJSPuufBpJH/DBrfXh0Dz3VhAaiOCcRC2PfK49c+
Vo+8hzaQORjxBfhQyxK4ULnGvH2/SW2JLQYBAl3QOYb9v7LtqNGSkkUZK3ORPP7/
gt8GjX2jNe0wmSAfw9bfrG4xGHNBu3w8HpdrQM/HYPDobRwXq99qy0YwG5jNP3xV
sbmFGPEHjSt0R0DXZ9oI0Ykl0bpQL2u90+VKmjJO7ABR6MLTu6U9vqb4HmMSNXFN
xBr4GNuaKFm4z3HFycEx/xrCyKN2wJszADB4dNPiX2N5iGW04pOuHHv0PqGm4ae+
Hu92TPq1EYsRRIfa4/N5EzT0eMY0fqNIA01kfrEwTUTfIeDKsXH0Ta4ggKKItKb7
eHiLPvHwJSAvXnPBwBpxqFbU9V14eBU7hkTErLhTKTlYSC0BZRQHi5PSugaVEDkY
k+nWz5gUDaya/eeToluSoO8limQVlnGaWoqDKj6Fg1utowOzAMU22N2ltmk8uZMS
Ag+Oh8x0lwXMg6EBgciWWQ==
`pragma protect end_protected
