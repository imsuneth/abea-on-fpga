// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:57 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sN6/ZZouZSbugOLnHdLqpW7M3lK1L+C1O+tbH9vH8N7HQ2702RKSRaFGgszM25OC
DJWkmQmPiJBe2WKV1104lkkSEHFy1geKOYeXMTgK27iqvfMP8oDbsNmzAhPE6uhn
/bxJlbnp32z5jcG9ic+jcbz4QVE/z2uGfsNZ8KbDkXk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8256)
2Q/WXJD6RAnhK9v6d6iqQDI3IswH+b11MUahaByUzp9tCEVw9SOQfRJyi2wTjhYh
pnae6wt0/n5GCTt8lIlPxd2WqUZgMd6s+Z9OnSaJFLNDkseYada/xSDgNx3QeBmV
yX8yX+DWs+majIdeACN5dLIfPO0fI2TRSN+1sHPFGlLdYS9cRx/Hb2tAShTFSSJL
n9TuxokDaO2ikZoq1oTwFAlppaewRvU4X9xWUovV7Z2k1nnsfOAvxYtcJxQV7vKe
+YlBPJut9/LeM/KOqDwGPsrS4m5u17TU0fm9Z1dyzTBhlalLqVk+U6DTyvQVRpL+
v8V1JcBll+5Hbdtm0r9tud/aMlkvXDJysB/zTza2RNxGlbwRY4TPuU+pS75xYf69
9aFdQ80fQTfTWarxM4/epYkI3nVlE1b0qI7QuxScSOZ0HGxCICbLO5BacIGBDgTE
FmA7JP4e6ypwzjZb5Ldqw6FKpnAg84e4zKrtPoW+ebqAkO/qlZP6pda45dgsuxlN
j1DJO8VGKMro7QEr3yJle8g4iXkfBtrJ3awkHywAWofua/lw4HUuwM/wBLlfc0b1
bIVh31zXLWsKtFTQfuMpL0Yq3MFFenZYyYC9+KS5SLaC117fD4M+pE2PgzKMC9uF
u/kFNtGt9P0YQ0rOQCvxww9A8nZIx1/c9f8Z0MkxcoMTj5QXyvUi/WYY4ec9PyAi
Ak7cmdrt4orfw76dNpqweiytb9bQuyHEYAve/9C182vX0AEyTxe5JUsc6fcTAlW9
HJMsU4r8/EVZbmmxXDtTA5EkoV5417qGrgSwdNHicgtwwtKiHlxuy2LSyNpwj+6r
wQcolKMG4iaw2Fm9IRobpDbRLIoTbMFPCGbOHDFLFzm9imNdMxxwTH+Qbd2Hl/Yy
kSop7w4/4r7vM9+SIjm26QcyxVS44ffwgGFv86/ONGJ+Odop48Tjq9ZXfhYoFj69
h7QCDsoeoid6AbMxg/qZAUoKkQHhb4EfalD+a85hO31LovZSBw7XKYEarIYWy8Ro
eTzKo3h7o0vTZVBkrYxtl+UHI805a9GMXJrQ9nlYdCSc1CA1IEeDXeB9foPk8GD9
kUTqo+HumrOHW4qmrqnevLSCOb5PkucnslkpCB1UHreKl+JLQMqXA4x2jbzqBnpV
jKlZBar9LV8saUsbXTuKIpp7QVGMeX36VLNOnMsc2T11ndByRscAf62S6eY8pKfV
BNFjiEuuX5XNkc24A8jXs0WDVxaA1L9U8QxQsh68sjr56fD1h4qZUoG+xWXc80Ht
PInNZuLlTAafi8uZJ7JY8+PwfKTP+gphusW/AKUamDePogHwgmOsl8bQx6jsH9lZ
CU4zRxusoDM4zOdaKtTplYlqt6QLOPP/Ul9A5SK0i6AkztR6b+BBb+nG5Dj9S+aq
j0qX5v6C/CgFPZbs5tOn9aEPiCLWorP/XJsYawwWJTKKWquAokIMYhoUJz/MLpYT
WlbkCtKSxFZ7fCFwjzja1h0yriD91e/dkf0Ygaij9rqDyKw1HZDUZQ3T+P7kb0QH
jIvKJz/7tH7g9jE/A2oEFhLYBg1W59IeUyrhxlMtetQo6jpAnFXBx8s83QVqcN5P
BHqM4W38TWQTi0UIT/CPJJmGy84KXa8au4WI8tlz1OjsiKyZaQGZR4eMhreY0KhP
H1U2ba10bZzaUZtVzuWJ/MRqMcJmBbuyHjHmAlaUarap9G1Ug4iQ+ddShG70L8lE
RkCg7e1elRcxJ1vu7B8hdfQRHubqmrFzWJCJYsr/0is+FR1dW7W3rbZ+9QJ2IAtt
isSL4ylihuRwmdkKemaq70PZ/PB4CBncvR1Yliu7qsRi41HCA4CZqmA3GN0ox0Tl
MeLAds5iF/WwPsRMmCQLJAdXUfzRL3yc4aGUGg3t7nbJ4Bgsn/dR3erjuT/2yGc/
kwCd1XSzxbCOygIBIwZT06NUTNPYBKFNxcEfdKLCWrI4n18zFrfS+AjQ4pF+Vc49
ANzl5xAUmLgTRo5E3BgoJumVea71LCvw+R65A4slrmWcjHrhhcq4oXJrsSI2RspP
Ni93fWVIvv2t5WmB9oCvrgBGnGySMOlJ9DJdTNJ3w/ne0m532XFhaZGEusrP4uqG
P3YehseGlERcJLum9DwrC6ECVxTQcfT7k8VDqIiBt1nnVuIpKa0mPT60pwQGsc7/
qVTPPLqLQnCXUfp1Bwae3r0FpyIoxCDCLeBfB60/1pjg6fKArxnF1Mbhj5yJorjU
MBLeL2espnjKOWBFJtWRYpJcA1ppR8P5HIQKZOQ1Gug7alwlwlVCSgliFXPY5Hou
U37HfB3kj5tef24t3xEuxUwoO+WwOONuoJi7IdMncNxoz60TWzxmDluNeIC+rfuP
vVlNYBefGQAP7kLKJ2hp9T/Zj7XqH1L2IAzr6i13bPDViyH6ktYyqm1XST3LshV+
gqBxsELpPnqXf92O0EGhS/cMHMZWcZ2jOErvhMWqdEGsZDI1atZiCAXpWmpIuoeu
qW4dJZXAO/AQkqhCr4xvEVMKJ5P8Tdd8UcuTYsqtXwXDA1XJf5O4p+8nW84are1P
mcV6hS8/b/wbf6+2Wcg/3UOqLrDbtuBEmbE4gB1cizPeOFjvufA5gLrzhXcJyPBc
DFgHyjyDw0wjddSyvNtOYy/yJULevVZfFibHpt93dxTHWGaZTPKrJ1Qq2pSS5l4S
MYhZw9T/fhmShhtzzRaAsMOe4C6V9SIjkRHYZ8gEKeGkBsfoEMvNUhyU5IzZ+aAH
Xk5nhlZDEXrqYCqmgWHT77qglcqhSEVzjlBprj6tlMqB6NOFCXuSkRMZ/umgs8Px
uqpFmMLY9nqVwXiCSiuocS5chTS09B3TJRC+qagvjpAN6G2M3HV2p3OJlVTuNNx6
8Nte3+crRPV4XaTk09/hoe4ci+fMsbISq5xmq89oOniwx8DE0MV5FGLTVE79fzvn
ZNkyM1HX9Ij9WkGU2iNgFfaFAYAiwl1sz8uj7PH7v/VFj0r3sJnh9SxIz/X08FkU
y1ymOENkvqaj85cxPKsgSgIOxL9poGUaRSlm3z3o4TwAyzEWfLr/cFVqEoDGX5Go
uPERcVUlnPgVIxWxv5j06Ff8gW7Lck9mKSIzRT2b+10VUX6y2VQHMQqE0Q7NCEAQ
M+plBapQlBAjOsaSmbiiVZtgQBdoukiMfVhQZCRF1gTjt+SKsfcqbFZ/RxbFherk
NRfi3isaiHap7E0tQWpoTF2b2uMXuhZR6cJr/41XBa4u/QuHtIVC3OcSdN1jlOox
jFv83r/y2aBLlolKN9SzLur9C8dE6XKk/Vo3sU2jT/dIMKCitAeUry9CnPvJwZPe
NroncP8ZXjvjVeXb5rmBbjmXbs8AaE73wO4SqJVgln1YEBwFSdOJmblzOgIouZ2f
Zg8rSZfdvcOuAo9Got4lbq+GRhDCGjzp1y65hCdWmXxIdzQHA07eGMi8Zh68uiy7
HcQccN4/rF4HlYWYK98CmcGPnxhyVByztB/fJLN4QfO9kYEQEa5EpV0n0IuEcSOc
6I1Xi2pk4rppXtMmWVhfjuThNZg2cA1Bqk7CmOd/IyRAyz4Ad443kbfLvcAOrKge
xCz0hD0dFdQu9FaNtYFre8S7eUOyDvjxnWJyUAlHsS0T8SJB4BqL14lJZrosJ/KV
xQn6TPwALXM6BhHgdKdczQTYCacyiYHaV3QP7hXzsYZkpGmFWDAOAHbQgONXhHCG
qSpZwMUIAmLe00mpi+akd/w0A6ZJ34LQ9nv52jCW+z9ytmKMsyceics8XcQJgN2b
XpuNDW+6/gUp40hNen+x/rQ1FrKtCYc+G2l/hj0L+3pN5ZX0J8YQJA8tQvn6LhNr
l66+HpQoJTTW3pWKkDVtrfPFuyNssZXjuLImOo4ewziyX866ziCyhKwqKQIyKNVW
DZ8S3yR8P+BqYi/nHqurD8/mnMJjQXs0yQhuWUmIMs6oqNExgEJToyWbUKMe3xnS
VhjCIWZwCP5R9tNILF9Cf1G1eb5de8m9kO9dXQufKFYDpOznLPw9RgIIIMRHknjp
/AkD56eT9iX4aSXt2lrwD/wqIJxCavan2mJ4kAW0s/CJatGpzht2vnRKNzBsBfsU
/FBeTkmigAehczEVeva6wsOGJknVRPcHcQARKQihRp042EFqMP8FjUHvSZv9R2Df
cW9wwQ8Si6DbEwHZUsYvNTWiYGt1af9PJVmw13Jklgyynz9wAKyk3vbzieebIuZR
TLb+ogCmYF3OniiOHpd5/00uAIJHsgdQsLeToByr3slsLIbMk2hcFd8j31iDzyn0
Mb3C2WQX9HGOccisuUeq5rVpj3PeBXlm0heig/tLQuPk7212v+boBqMWQ2Wm25Rw
uDAcxvL7GJFtqgmhkbTMOAB7f7bPm8tH4x+leGEb0XxRFxDvmsdd5sQnJikgYgcE
37FjJvaEGr+K6Umh7PlpeKRBrfBnRZDT29lzDTSzUVcN/aXYbWKOQeDDoe+4WBqR
mFsf+nsxvew2YerhoZs9G4Tht++E9H1V8IUsunsAgZsTfeiSuGYRnnfhwCYWdpCb
IuVW+qXT6UWnKO7UBLbuF8N2NRyeIPeBvYCJauWgUnEA2+lsMECS3TCqedEBHrec
Efr/K2EWu9KInCZq8RpIb+hdginWlJ+zaNU8SBkvKTx5lxdXpeq+0L11nawzJXeh
yL1x0Nb793JRAp+EfyY1Viewqf5giEtUS1mhRkU2R77q8sntjH++/EG+hW2SHPMv
16W8a+ZepquAv/Dqu3oHoXZRHhX5EPCkjeEWlcKbMiPEvPRD24PhrC5BWUFxbq7U
cYztZ3OvPNGEYN1YgDTZNzWRi3h2z43t9hj/YVAmDpM9s2g5IUJTaeXKGzVnsdBT
wdLgnlmu9bzADaO4a9+zFqbBpaZOIj0Gv4/TBdWQrVUi+2oitKo8mijHOd592gj6
bu2Lj0PnI6qs8Gwl9/gfY8zRp2mltQgZ/hQwG+OlZW4q3lQms8rAIynjHxN3iQm6
L0lTjIT5zIHHP28L5+MLNvkOhejIgQkfvbRBaNKXklJgi7Frp+w9AdKes+UXhkhC
dpCXisN/UTGh210WNploKZ50XSM+Vjz/h9Dhs1X6NUNMdwjqCUh7TINqPuBiDSVX
Sl1RWoyy4qpvUo0Xx78knvyF8Bo2iqnQTWWqdTZqyuJdfpjC4wShuMMDIznWYl0k
K8HhNMC7G7eCZ4AneldNm5dXjfG72IXcSBflMVE4InzDLYqlDfek8KILGxFZg5V/
YhoMCVvxzto3pgAl1VJsz+BAXFWn3pAwq2mtibiSl8kXe0LqvvZSb/pyWeXO/Nlb
gDcGDoLcKdI5dFWRhkClrnWvofAzMkeRJHKavZaxExLxxvqPXP1n8nUZHs3UUlT0
tgDw/ScBTA9bOs53/qSw5Zu/nOiSvx00oQWweIDq8H/kRi99hbS8H9mlLU9WL72K
MLI18ueO1zk/0AwD01CvcurV6BY8SvMM/vmDUqPze9zucd0dOzA9D3y7Bn8sK5F1
KYsQawuhi4kd/SevEoaWayWdvxN5LwGzDjQiqIJK1YRZDTyBKFTlKDUI/6DKq0mC
jCji9ho6kEW0dIz3q7UF9zWv+42N9ghFxqBsakiB1eYcU7KXMOfafB+w1F96zLCO
Ne7gijFTLj/xW0+MNZRVoBUaGIw7eQSsaAcN53B9KJ5iZZKE+jr/jmUUw558ab/j
cVelVLHzGIGvvbrTr7vZsrUvOXzKVYBpknU6zsLMu2DbHruuh/JsnOraOy3eLlPI
93gYr7vs+dUrBT4tNTzmFYBuN5rfJixlM/nwcTtgI1xh/HVKq7Fv0rPJoPnMqYm3
WXG2VshS3Y/kdWwWMhrQS+HHKHAJbKaFcgoAy+6V7OSQIFcqz9v+GNFuFxquhEEX
MUSVZFAeewP8fOkDDCLrC4EW535AIZf5+5ywrwuqQ5YkXgzkbIgcapKWrHAn21Gb
BcCpgabjZWdfIDpRT3V68KQmsgnp0JFzrm48ridD76bvshSzn5BjhZ0Mgf2mE9Vz
7wpU5uU5pqe353RKwjMCFj7+4Yv/8fJX2l/t4nWRXnV/y8bNJpYBNArK6z9ebLDO
WcZ/4Kv9CqvI/+m74CDug6Qitb0WAlMUdy1Bs6RLtoA8qzF8eKwIdguyaM2SyZWL
qhZU83ysxFz933KHYO7FuK9OMM5YF8HpEzY0t5Fa1L2DpkCWz2owF7Uhb1j8rVdT
UwJfA5+vSY+Gh7WH66abBBYBcOp45RKeRAGuEdgB6Z+vkd4YCOQcLcmfyJxg9m/k
uRR7S0a76cyGNE2KMUMvGZJtoBeAgE+CzAi1lZyYbguxAKXy+Z8ICQa4002q5zBd
CVV9s8TUkOb8VHGL63UrYE4ZzHAHQcBIddMIN+Srnlw0egfv3ZqOtRTdmkgI6R/+
Sp8IaTyyD//dniCuN6DHzECdg7UVpzHPBzGpUya69kU4GTBbnpJDJc88D754sc5x
QzW3febK4B3BvuIA/mteVfkrttx7O9qOjgKa0drX90A9IQMHeWgkLY+C3XP1WBFm
oxJB2L4yow4/CB3ls08UifyOvsPuH5tyhd7ymIS8PDwbiEGKFfTPBCnw0C44JSKH
CT8UkCIr3tD9yVt9J0hiKcNbDtOeT2fZ5VuFnk3N+zLYTrWJFYbYDL79Hzc62Rsi
rY12UEqFL4Xm2yB9IdGZYmuOkFl1eEbJI6qdfN8cUSSM0a0ki0eQNBUu7VGEU5cJ
JVChMbAcKxj6pED8iC5O1gB9v0TYA4SZmwlUgY+AbvRcwaAi6zInZTE1lJgLx2mZ
JVEGLkQF0aWtH8zNMKcDYFSPlp2vfVsNseNZm47sidap9KCbdVIC+0FefZZEzyIq
Dy7nnTPQNq+aGKOVUzeFHLymAxhxHAPkffijJUDZXl35CICRsOjJ97gxp0UiJr9L
Ftn9H/sSveAPMMLHV0ThLZbq3CJQD/Efcgt8p6zEX8XkWA+/4s5MTNn12X0/38JB
yLyvHoBVLRfr+z7ew0h7Rb15miSUc3QEr1dtkBW8owb9/+Pt0GFZhQc99SMRDObe
+HRDP8rnFRnEgNfmBQAuWtdwxUYEth/PfrZWvFcJtpNnfJ4bkENEzwlhSDLXTznq
t6ZKiN2Fl6/+20p4tZrhMKwhHcnBcCtwBywYxda2MCybScDRkG8HyU398q07Z7xb
30XQVisikmrZCAI8ggm2Pr/gon6mvZkIXMfTIUXx+AAOGTwLBE9OmJgO2ocP24RS
Ho6pk6nuFAjoV5weepE6ekVrancA6jFfJizOgsGwBVp2g9NL/5Z60EUhUGJG6xhc
AV+AL4LUCwMlR+2UT2Xl/+uj/1MkasD+0EI4KBMfYY91OEYE/HkhgPCSBa7pfkT3
feU26blqfCumXWmnoLK9SQ8ei763UF3D7W/9KlJEaQVH1aTYsrUlw3IH3tYqwkT2
A5LN50sXBXihMDVTbDIGm04NZX31lfoXxVXfNPFE7YbLud8dAhCck+i2J+ifIRLv
tzfcIfc27jqn0qKjdFnnzQJpRPfbF/rtFaNMjYQEW3NTaheSsQHM4JVz/02SPZPz
V2egpP6Lc9kT8lahqbvjuVPYqSY7DeuZuU9Xh2NjRJTkfVAbaiAvXqnx3ZYZbNnf
epoNCRYq6FEeaL6cWsHyy6FQcGDhdj0ste3O0h1yXipdtdmYlV/ipDARFC+YIkNR
zVc7P2Jtyuuk9lKGHBJ51GT0D6OXX4hJKRObB51PqSc+e82HKJ6/bFDkxSHjPffb
Qc5bmx4k9CxPOO9qR5VrbIR/K0pvc3gk3zTDmqSebXrH1953e1tYbN9S8vykbX8A
g0KiYXZN1LP5bGCqwcc3I4nzw6moLVdZzQ5rVE64gdZcYWsUPFHvOnUpsVTsuytg
YSb2JBqVvLhboOiPg3WOY1NlREq1LyQ+NqbTWKY+u867qfVM30qq20XP8EhtHNQG
FGkYUrYbfj0tlA+0twFE86C2UbdvWAeollQboTnxhhamA6IepX4glVL4oAmVWQf+
h2sKIXMKnX4RtOTFxYD5ijFica6gt3tinPjBNN3bV3hfY7es7zSzfeZcyV6rxpby
cL1xrDDED/G8KHnYiCZK3kfwLNx6crENhx1mR81TX5gjI01hoJFsf5qeszEYiRKs
oEG3qzMJ+UM6P7exCr90nuAHymi7PuEFT5IoJnyWxxM52GB3MBUvVEUso2xSLtPR
7RaXJBb0GaDvsdyjYc4iXjfQwqkqsZUjWqRTvMW394xxPRKLsu+m00t/6zrDVtf5
45dlD+iLEKoDLjt5kPzhfKH+803SgRdLgWzBxiNSftqAy4wAIC4UGoyMRNHH0tZZ
AiD6TOLvWsQfnyg95SCqKbk6g5DvUDQxTI0ocxXcpoRzGl3xXkxr/VlqiSptt1JV
OIieosfjW/OJWOEumLkC1ZgEurz1BRpMcrlhqKep4SxACO0f9SoIH6KgU0+KWRwz
Bc+NSEZLnHx1TV6a/nic9ACGnx+cADe/n4wdA/XEDBxIgU2Har5qSBDPnpzqUylX
45g4M5i/IAsSzsxAin6t58N7O7v4Vo9/ogCjizUJXdgyCBpk3c6feh/pcf8x0o++
fx25rDNR4NYf8t4kvj1IkFaai44dYGVixsvo0eJhkfIH7GPQ0VLEpyIHg+warP5j
1QEOm3WF4IBedPGwcwBP9F+E/nL5aPeYV92gZTTGyLi791Eq6v+5RNkqGatNAwDl
7W+yUr+d9c5ON6W7TThhUGzHJO5fJSubxXHRZfa6BRuBP0VFdK+uIQCQbd/FLgzz
osjs1F/f2LlE1maOrMh9HlPJ0WodIEyCKPR3PnCbru5jawtql9Jbb7+XILtmlbQU
2PwnomGHMmkLdG9FlxMlkYUE17CMf/2VFIei3AFWh0AB2BhceB/bL5RE94g3RnEI
WXeV8HW2GAESZb/FA4MxoEv0935SXgEDOYfWaNU5r44BGuzDNE5ilsbXqrYrBSf4
STh/OaSYvV2d0x4PjVoKwJa220bB63G7vOBpfALx2+6vUZAoKYyf7K4tTcHjjqtm
dU50u3jbduEfKvrccgSuulP5GgR9ByTfgIDqrHoU/EtcRudLBU2dzaHfOoMlqjMY
uZLxT2e+O0cQ5BkjGrjPl+L4oWTpWA/Buf1q8C4TeqkFT/I6HavYvy/pKBVyFzcs
VYyZkZoRyOkidczt+Q3EEW32emlI+kMekHC40TotJjh80TpVo7inkvhsBpMnLiMc
64wgA6xBm+soCT891vxBtFjuAJMAGy98wbKymnjYFNCdRc0z1pmCbBjQ3a8zDRgQ
mxSj61xa+Jj2+Mv/wvAWBsnkx32W/UPaWmhTM/m65I26b8/HQhZaOO7qCFj9oZp7
PC7NEpfoh4WB4hy0Ofp0VNtgVsqpI/YJ4rcH64j4j2RejqCQz0Tr5XipA5el30cn
4NMDQuaRU91PQacfQdGIcrXV0aB02J+FHABmR1U+7MWCY5oznLO0Vy60Upq3aOfH
W3oromyhgT7OqmmeVKv7yaGa1naypnaAk8mOnC7IsMtTsNJViTMtrWMKLa2TId1W
6BPTzNeObchEvNZ0mgYTD044L0Y+Au5r15cB0rVfmFfQmx60FYz7gw2YMjvO48D9
Vc5+b1iUkT1W4DTCON1tvGsQltXFY6Qu+WosAUcxtTZ6GRIvdUBBMgdtKydXWUyH
bQ5R7vd29Mo2OXFU5gnYDCrJ4uM2+H5KJhnY2K5JxgWt01xwdyV6dqV4IL5Mk7l6
yNbFL/fEsMHaGrbwC/38Q0MuTxpvSINTm3mbzC5dBnNG7D8Vq2y+LOKcYjyhcmvR
ib2S9fsJ3QSShovujiSgqKlIWy9fAI2+7cjKDSoRsgvOfdIdS5mn4ngod0gv0xhV
6I6SEsJ6Al2FRuVNWT/uazz9K0KVvyNoW3M7Mq//ZYeQ1RkMjHbnr8Fz6r81dsab
sloFIap/0l5afEcwpMO3p7azh56m0lYnfw3Et6szExYvduhTp6w0K3La7sj8NG0W
dwq6bAt8jY1RPjEQ2NcSwGsHXDCfypwJnkpunBU17IoZ9wDJWoJq+jAJJ/iwZYEv
piQyNoITZebReyyTNSoI/yh+zJzUtFV+CyOkFLW33r+tlTLQo2rJumcgoJhpfVEa
pKjmYvMhYtatC7SquHJAxpfPM7V+i9joROFYMcm63+0XiQm+ijBZsdtxFvl+91AA
cHXHJ5UPJrx9lNSr2hQQkCnZ6oeHVUbWiFWJBe/8PBFeKHsl2ZwGh0xNeMf/1TxU
VGHTJIpfpJTA1Y+lscQN7+J8rrH+XM3r5gdouAswu4JsFbMkwnkEXwg2vxOaQgYG
3fD1h5ymqLnsFj/DX/+HSZDOoIuifmKJXGSpQvmJ2OjeWuEzxseNxZ5y9fy7aB/m
KaEF+uUBXajJBce3+nHBxYtjNSLztjrGTqDYR3ZBovGuwFF3ghUVADr3hecqPvdI
UCj5fFhENZRIa5OLhwf0kVpvIIHhtZ/PvAJ+XGDcp3z/bOEVEndE6P9ZL5VW7h0e
nyNLYU4OXPqwIHC67pWABEiwgu8gjC6JqiUZAG5JSwuly4jrkfxyLu6em81Kk7mJ
tfU13oOQZAtoP5mTwTjM3HE2/Dog/ZDCysfu8BzeijhC6Psvj3369UYxZYqAwtBO
XuOC5pEpmaebeG8FxF58ledP8p48bNU2dB+zVWgsKrvGGf1fAy8mNnomb9cstnmD
1PZFJWAhNVPUrarX2aVxfws+sDwoLl+gyTuiaGdYnhHkGsjFrF4nnsmeRDMtFYlB
Qyl7HHWBQlrjaVlYw0pkZ2QpIXzTEbbw73lDRwBlzTxc+pOr8NcqvAkLuoAzhdd0
zV0TzRGshvdmpy85FBE45YHIWtjz3y/+ji5N81ljVQ102N1U+WpW8sO8N/06SBGc
nPekcC4xrJYyi9PVQX46KgNSkEQYCHvZypwhEE6RuNdq7al9EQYPvZYb3h1sK7wu
U1XdeiuPD3d8Yjurpy3OCq75uvMWGDftRX75SXdJuf+cdwnDRzroHBhGt+HfTbjT
`pragma protect end_protected
