// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HRaKpzhQeZYFWT0S4sJlDNLo97FpLhoN4DzSe4KIwClO3iXdfp/57gKET0GN7lis
ojMQ6Gsej/en98eRbkiSRqo+adPDCZZwOXZv3NKQyKnVH/outVdMKYtxY9SPaYRf
np064bIiPbujF0fYIvSw5KvCL0BdX+5B68aFSRpW2+0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
fkGT8AbAovoAI4EQ7BpOrgJBFJ2donsFGDu8K1MbXGKXZwxDBUU2kWcdV9GHPkNJ
aCgfqc/FoRZrKxSB1GMJuF43Ehf59XsBPc7pauAfT6hNu2E4JZjejtw/Mqxjgex+
UqKqojzGv07mMyrkqCcpvLar6g4OXk9KQlB5iL3Gj0EISxPHmAqcnyO+VhCyH5AF
ZCPjXyPc12fXXkviCUR6ngoooiV+etU49iKUnEz1uq3AdZjATMm3XG/wLonDmPGf
ny2tajTFXXFLHvFQadzwt9MkfOxZtFQchQXIm+0lxOVHe77O3F/zoajZV6U4/9VP
7tvgZueLv4nnCL8nCJKJyiNsDRXvxrwxHKAVAq+eXWavJAq1bi9KwqQqYMYy4kTb
IBWdsXbnNHfFI9+D+kRVOo+6SxKs6lY9dFpnTLwU8kbcUzMDcdVPJKOjl6wizCX6
WWt88wfbEhOQbOFmQnepm1Kd94uOwS5z6xsqtH/K9Gdtt4d7af4Bev8al0O6S3Z3
dnk9WSRlV59/OWt0RLj+nZO+OUb5AGJ2Gbeegz+dfCGySnzuOHoivLvHCTCpk4Fg
41h/1pR7GfPwwanb5C/aRA1DwBmv4tzLAVOzQssm2pPTcWlFBVJfQeob59dUMCtJ
bCTOwuffDreLuSqVhvfnrnYf9K6/UFZX4QHk6ANnY0ea6SJINdH1vZiKg7A2JCSS
EcGRlX64tLl9ysGAPM8VIEljFTTcRLZ3QNAAKWQwJuBWF4isynmvdCOWzMT7lv/d
DtdorvNv9XPwEUcfN0aJvSmsJEQIjZb3VMEeHl8+3qmVwdwUXTVSBviiX82NU+Vw
w2G1Sjkcu6WyQDihluvOdegdIjxxjviJBcgVBc2UufKoGnH0lOAATB7+VFeJwVM1
ZTGST7takUo6ZxH3VxFFnXA+1YjbVoKPEAkPIu59PzlAb3hUgrozEztQsYQdXgTH
/2AiRCiJGB4m4eoXsIhsiRytR+wjdaIXhlokDh22NiSFgU5UZaVTi+8iZ9T4SSya
Tk/JtfoU1/JqsnlqdihPn/C60nFiXYalpxDmeJS5e8/KZE3JEbKuTo2g5ennP1TK
wU1mfOzGi4bPLR914r3IKhDxxowubP7T56B/xN20bhcqKs15YIJFwlGDlYr+qnpk
kLf9ozBTNIyY+V4aMnu09MXqGPzdGW+JWb3iZ9cV9o92Y7erPpSK0FLWaa2X5iac
+9BwIcwOjxr1RjBI+5uEPHXBQ5D7MlEX+V+Hq/WRW2Bjw3CNjAjlsnfo1hy1jcdv
7vVSbLqLBKIBgUpuobEaEOzQOmGdUidSp/9Cl0SjY9UfWea6mUTkXEwsPeMPgvMo
yxBxYDY/n1w7ygSuI20g4Ug70qkXvM08PozI7BGyVM3YaInRJ3fSnASx5chxschz
SKeaz3QXDemgkgp861rKkEpH3cIny4Lesnw8BDPaKozddsikE9xHXN3u1WTL2sYw
HO/Q4kXkJwGaKJVM4YjUJ0IQWbikfrtzx6WE0pipmgME//k9IE/3s1N5Xku66xKE
apQTi0ETMXFfIKhG7hWj/9lLjsaKb4cGVwfmpPu59EwhomCPd9XnYwn9AAiZdxiW
sUZRb4ghp1H51l5M7jwdide36E7P75VJX2Wyn/knk7moyw/anm4uvSxOoPE8tyXP
n9qWW0UZH44n17I0mqagyqUnrknrv/Yv2qO/pGGPqQlobk8HQjCwR9fEJ7615zO+
yay7SOryskY6rugiFdSZFsT7r/4T2/1B3Ao9jigm8mUz8OtCV1GVOd0kwctqKXsW
95UafCxD0F+BNjG9jhNDr0w1+HmgVO4cZBzkklRQ2cX/+MK/OrebWflEkKYzsCc2
GzICeXreRbQfEOwI/bqZRGtnm5jus8PGbPuGrQNg6yvEcsXnCwato6hWFUVSsLvU
9njpZa8RwXMzp3dwd81tumJM/paMMtjGVPbBGYMH81mrNRRMUtNuyVPkmzla2avM
3kIno1Ssju53++nG8RYTpT4sbIIc6e45cUyLTW0FtTwWiUcoKLMalVdkD4m+T5VS
+z6TBD2mpFIY0nAYo4tfHQF6j2ScHRjwTxA2kUHlWznBZ2Er0pljHobWrf7bpU7e
PPniuiAFonmaFv5lAzlMB8yMQe7gZyAbXd+v/QjN+Q/owQ+4vwiwhMad+FInd7Ui
XTdCXwPJ+eKa6uIEhqp4AgYWN9WcfYhpJZbYfRzK/JKl3e+isB6TceRfU/uyd9qN
8WwenwPC5212dijea3430rHh3QWNQV8hIspYy9SK77xOBdpBlRxQBjTygoHSfnnJ
nQtuX+wiIhOj0oJJyip+puc2CdGdDcsAT8nsAZQqkQWvdLF2qiYNn2OAf5yEjRx5
3XogvZuyioM3ZvUVePUFAPUKxpBVJ8afTIEI9uRkHmi2ALqjQXX6/GzDZ7TIK0Lw
Idxw5tukfmPcjU4REcsxszjazRgWD0SS4TatmqU8ZefFK2JIuiyiew29FPdGNLAg
e+H7YGeX+Vc9FL9DlU1OuCaXyCEU+VrmDSXc76qtjxf54A7bIUv9vk/TZTjsRUjh
3pXyWMxw2dsehoggG825rUxzd2EmSzhCGGZIu/0ekrNPM8g+cASbS6VM4VEzl8Sg
5rXzDT64FvOVmmgkQU0PjfZ0kRm4o6V5rKLR0Ia2Ttqx2TmrF2wTwGPkrCzLcBQG
nbN/CLa0KzycK29uEYoTDH2U0G9UjA0txMlZGfb0M4czLZLuojWdgL8oVf2nR8d7
uzwTeUvQGa+prkAQoCK5bmAU0IlP0Y41ujUqYQFL6kOquruZQ4Y4TsUCKZ4LJ1UU
jxuXksWAm2g3SGlRAyJLYGR6loM4CvTSqzd1elYVisWksane5uQMEfFqVyrWkfJ9
IoEz2tAQoqxNuf/7/shNiYHWrgmsa6Q9/vHGhtyo3P6x+E+2BNj+4nS4G/aMynMZ
M1i4oivVQAsEel0U+Fenj7N2/DXE6otTb2zcrh3PiRTCXY6KfcdxV7N0FkjFl9UB
YSfVI2CQQR6kUYpvbPuVbXoWx54/rIZsSloan7rGZllLFKSs4ESzhDnc6SxjZuWs
FdC1P7LoisfJttTuxQHdFLvlvTDcA896U5PIl7Bgy8gCnfwUvVOsUnF52B4oZuu8
q9cMhyl3CmkEUCZFLonLG9pV2OvIPFjhxfrzG9cFFXmVGM8NHufX0gJXBOrm5APW
4wppUWD2exnqOtXYG0l7Uv39EfI+EaBbcw9f3SfZd7IGfye+CDN4zgPQYNUuxEzv
ADarnzeaLlbR9mUzov2NWkwhHn4Fbwe+HpRyqr8zT1+AYyXNa03kaTupHRwzWSiu
Ao2AKVifaW4yoE2nFXl1GpFJQnXDuinOezixnA+3JUGaPOdmLj7HN5lHQ9GAZhVY
OqYgSHGo0tjMxExLmgNJEc3E8m6SjLu9O3jVHS9FVvRwThHBZ5FOPHCPu6CIrnJH
VTfyQMRytWIsrbExQaIDEU5GuyYvz+c3Sh0IPbo/Ff92mUA/B/lgcrHRFroTexTg
uIZcQNDDD77Id4Nuix3aJ5dBMyu67BdokCjUWF+ANzCqs+rBvbtwH0f/u96rYxQw
V7IHR6ErucZSP+I2Qwn6LGDLR+EOSD4cD5Jth2IPmOe3YvvXsxJeQfKnMMSjXjTG
2YBPhTyFQW/CT0jWB0ZNbxJLerBy9VOaTYrFoDggxG9Ki90Ny69Rci+uGBKupFlm
ZAV39vO6K535hmJKkqlAlIZcpEhD1CVjnsDhv/eGIRAl2Os5G+UrgkcZ/tjmxp+x
IGNB3Gkya/RrpHm4WJsioxK2pdCDYj2ZjO4yh/8iWq2nhhWU7b+ZL80swKpAC666
fna3nblyRhWcnK9O5OePJfe0qdM67OE30RVnXWd7Y4pGWWUn2qo5m2zzbEXYvZAW
6oyiNKjLvvoSKmqeTgE7lhLtwstCGxcFtcJ0GQyi6E0mJojKEouE7ksTIQ8AjSdU
d6vjSjuJbzy4xz+L/9WvvimY+OhxZ+wYzL9T6MLqsxAKhKOfDwAueN9rQwVbq5Dv
BOGUonBWhxpGI/Ofu8r22R93jBl+ZviidVMtBWHCkM3VdJaWvsDL6Dq072ckYczH
kwPTRaL9IoOXy8UNaXbeFlbryQwI6mauNBJCjv3odzA/5nKa+8jzB+TeffKPqwEo
sSxR4rRgnbT2kw8bq9s9sYHr8+QfkB8qQzxWIacI4GLlR5F5X6u/XKcIxv7z0NvX
7i4N07SKWq9S4Rviuf5iCssCcdVwq/hwnlzqwd7hG7/Go41z/Vv44IgzHKd9b6P8
TVJbZnXlXekmKUgSgRzhszF+2VrPFarPz7cL+nyLLz9qwD/vC2fziEkh/dUtea1g
QrX/RfLWkOgSo/DPIqvNlXxlxbXQXWzTWtYDWiLGJL4duYeGnKLuZjeRww7e5Yd7
jN7VDauYTKy6MkGjqlYX8Sigtw3W7SMWtlMFZ4QYbMngKmWo43p+Vv2wy7RJ8KmS
C8q5T73gLx0aFkfHrOcomA6Q3nTLOrZKjZzfQEAwqz745cQ4/FxuhCRhDDrEyo6Y
prJFOntFaBckJfhjHx2/vIegYssrx5al6oxeA19ODqQATOzLOhYH+0DId6OcFzDL
HQN0bXfQTovmNz+P6WFVKZE3w4Jl0IoZJS4reZYy3A2U/u7zMrL7kxTcaI3XKd/E
6I+iP8SB2rL2LFxZkBDQMxqjisUWNamb/Hb77U1NxrTTC268+y56pIRx35flJKwf
fi8Jk+mEXTpCT0Rwij8spC6vXudwaK62dxIiGuMIsfKZfmU/FVUrN3Rl2Jf/JEhs
R2rlhOahN16uXXFYTD/GtD0hMudU40MXs6weKueCZba3VtWmi6HQPhUGJZuGEQ19
8C6+XBeKpV8X+8fkSpJFfwU7x8PV1wI80HKFMzAw6QO3quTSEc32YjNmAN2/ZDn2
vAjqwwNNkUJSTh0hfEMcO51etMvNmGAWLAr/3YWHv45ePQDsZQpzM/nnRJRfi1wy
fq0TNAPJ5HIS6/NoZ2+u5xWtGgSommMCQ5Ayolvyun0KByUzw/E+cJCo7676hL7w
LZ/+bG8U4IuA93O09WY9m0ggJ/8Hhywit61MNz36y0nMeOGzRMuw+C0Qd5jmhBsl
VNqZLkNceT1d9FQIgF4/47LVze/oME8o6eL6l2JS4rWwkgInhvOoSXLpxBjxPsm/
w0UCkQ8WzPiygLPa0f68wNkx67TtmzbjwdZ6AnjaureCB2LvDE46P9MkmGZUBvIQ
WGN5J/PnCo57dyVcYr002RkeMUIewpqAmKi1I/Wb2VmbFwhYRehYeAG9xchjPmRn
QI6VVUnG8nyTyH4SzEYbboj+ui9tt+Bylsy83WEIzUIVSi3aieZHvlyvU9226c+f
0vfP38uIggWEqc8QWKuds0QzPfWxFAhdCugPVshqcADouZGt+Gc3Jhhc5depxzcq
NC5+GV/X9BCOfrJK5rvJG87B2GFin8Ef14YfKl605VyCHwOmeN4Q1x27yQ+vNaVB
qRbkw908PFe7gaN+y5c6ySFmX2Tqe0TPI/zrHluqHIic1wK5Qgc1gYlFD38mCOC8
3CyihM1nCPbNYaDRLVNdyqvNnHy8X48z0FsKy/eFMUiSZ96nCa/cSvE/cNNoZ3jB
KHugr9wmCoZ4VFqdVUtbUC9xGADvWe4bk7OqXSUw5BPlL58ADLEHts/qoodCaYLK
omjcS6B7/l750MZ4p24uTPgpUVGeXtIVAoz/ryuuZCIWxxBvYw1znw4/B9CKxaK/
kNb+yDRWf6K3IUzevcZNg4NaV3T32F8i948daBS4TxkTk0Y0iO5Z41VqdyQUIruu
Yxx0UUT3wYPSv9r3iqJehlwUh+tbjknndT9N9JS8ldwQoSjauRT8cezhv3HtRyP/
Df3c7bAkFYxkkz0uvmIumAoargH4e5E7yIAp66Ylx+jZMeqe9PYx5VZvF8nNEQ3v
iX+PwCTa4a3gvFVdWtPMmh3ygiMvoC1PehKZnbOVD+Ifc8DYhAtiyxYwlDoPX9tc
A9+AxPvABnlR53gfsJ7eqq4yHUZ/MwXnysJbHAO3ZPpxN5snjItD4uetDzHcmDI7
yfMM/WpAKAQ8pyQ+lgiTSFNXXGBzqEIEj87nwrwW10Spg/RmewXdMvG9zvqiyGOj
C6sKJ7qIYbnqHhRUS2nTGeP8woRVchO3FGbApIGqA7Ed32ABe/f9GDSXgptqGJVb
QMDrJg6RKRWvSS8/dMUwhfxKqUq8Z+tT3OtHwf//bGpJ3jCXn7ozMVJfAyrHOnHS
jxcTao/Cj3L6DNU9nwA+nAfCSuA4LE8L+7bn7YG7ZqMtFGe3UdXne5FLZ2QJkoMQ
jd/cKxORoYOfy4Szt47jYtJ5P3g3XiSJMbnRgMCHYnW/UYnJ5icknVFLWN5mtXcf
fnq0Dmh+dOFFTpkhmLZBMq/tEj1Vd1Riep3E7A9/dnTCBzxAk05YUzIwOIZj3XLV
FJ8wWfOxHU5PLiiyJe5lt7GLpm9RV9Gw43fiWEM+ALwWyIPdZF5dcPt1P0/G5O2s
XGQXwrZTHZetKj/wutMi+iwVJPWXLgH+HgjyFdoFqDyMAycmC0tyxP+wzg1mZVvF
KI7xcAaLu0CfUi4Hov1eojooRYdGfA4TTAcCftZGprKZ1OvvJR0bSnGCRzz6atx0
gJ+6n9kkHLetqhobxed4DrblDbv4ju0FZSnc4/dPnbH6lRTnDZ72gKzERHfvkN0R
M8ZapTZKi+SpqzKH6fBjXN5YDo5nyscjDFAtVasLI3n79eOqlzabodUaDuePoJxl
6TjDdmN9z3ZrJ0Q5F2dq5l1D8hYF5yHFd8k+IMxcdhacOHFWALrlfRJMIX3pWfj9
mlA7v6bEVEVAJvFsyGHDqO1jl/JVLGdRoVIft8mcD/Dwdc/XmNJy1N92uNYCaoYM
NvVRX3waQRuBQKFmijjspPydEDZkLFktlrODIPKFbcAr/E2pg5UfM0j7H0QyuJQf
zpYtd2TqVivet8vjVWYd6Yqi8TGanA+6HS0t3G3PAAMqbPCMFqJ6AzlSLstUM06c
2IGkDTBV0pkOYJYxOb+FlOYh8W2vQQ2XCr6run1ExnhGr0v81CCiqWTq/wlD4ixk
QUvUF6VBfxKeQcp5NrwZOW1YtvuL/51BiwI+8euYmynaKIyifqj0EXr9pvs9ZqC9
Rs/MX1kFUGIWEzTSgRlVFjzJsn6srZSXGIVPGp75L/njE7UQX2ygnAQjjMB7BgFs
PrSUMt01iwiKfJSRFyEY2wF/CZCiQf5cIDNvSx4uRKiIzkxUcMZc9a4eMp6jgzXk
gN3bV6FN+x4XLJb1mV9JFx8L61zGKD4vvKDiCm0kUheLoAcMBSwvvfMtJErByRgI
hwoR+3ZGRNYtwR5Jo4fOzfz86ORARf5wHSTZ3/v1832hmpIPvsR3legMyXHCcR/B
pwm/HYw7jvV7K485Nba6F+q/qq/Nwe9PEtnCFR3hh5S3zcrhGJ8XI4Cr5VdxEwll
oJsHrQFXBM6d94sn+k38DCGTFuI2vvIWEPpFGE4OiuoRGDc6hwXS3PFwGOH7oOEj
fMLrVw+ssg/+9rhixk5hHHOUUE/a8fXX04v+JEUHncCHSWeR3916FmybkrmYv8A3
cfDwiIk3ne0GbWR4UU6PUYRvv/Kl51xq0Cgk1fnRDJIpXr7W8lkOJuwIldtDtGLO
Xda+P8D1mvmXubimpidzPgTixuWFnL3pAMw61uwUQ+bYPSiqwZVhxnYjKxq0DOv8
laKp7SOqUQyd4ZbVronUroHcmujCPVWromPbw+7E12KAF91O4eb1tb5yZ3RlNPK/
8Gg+Cmm49CZHVMBi9CsFku+dMIMqWddzRoNbxwyeilAIYEOcD5veMLRMLGvHI9x3
l/LLwaf4M2F5FC47SkfilhAn91U+Igo3kNmD5nt5GpxDklCkNb59Xo8aTgNbyfya
iWrCFckL47Ogh7VkqHDiX70UVjbL+gw7XGRRXzolXUaA0MA8IidKUeoctIkd6t/b
5NV0VudFIxxX/VOYxanL1/oulbSE9I7hxDN3khrM4TBDDXwKExAJr7960d/2jMIo
dHy5Fq9CynqOzS+qtH16vsZs4Yp7uEQ/VWP43U3/EeqLKGh+byg5WVte+guJyhAf
vCDXoCtXQzyeqw0YzoCOKe0A9tgLhFrbXh42gJifxqcz18gM5KYCU4UuInccAdW+
Bl+EQwh6F70+Gt38ROpgU7pJEIhz55HD2bzbS0ke3f5xFclyg7naLdlqOJaJaKDt
A+aNzdbm5Vy7r+J6V4gaAkwv0AobT5QUxtp0AyUfvPOH7RpoBieh9iBqcFgTUu5v
7zpNJVwLmzooiFcnXL0ilUAeJjlylNknQqDuyeqVGLBjDZ03F6oFa/7lM7Z0ubt6
xSHouExJTvH0OxHj69am3GsdM3tks/YkDksIh7bCglKFljx6QvW+px0yW/ec96Z/
WHOZI82x+JemU5WIvnoraTjMAE+uC15z10NQmZg7YC8wtuAluIDfSOLnK570IU/k
AfPrGiUj5XlTkQK/FfUqNpNLhBEO5WyAgWqzcPjXc5QywWyrnrykWYqynKpeZA2H
gJbr7hXikk3Aal6yIJBixq62ws+Nh77EtinaFJc8+PzA4aaibS2wOdBmVq1+TlBc
GkUhRMQGkg8jaWKhuWDfHmnCbksiTI7wxveIQ6YgTOYlnO//yzASIwwiaYfSF6BG
4f0+I/v1dML0eQjEedjEreVCTphtp6B/Wyve5QPQuFhm7ZauVTBUf9rDfxQk0ais
uqqplakphz7nxnoEwLdhQhSojg4qUdBXn2nFB9u5cyKN7nL7kYyBZskVuhSkNuT2
9ZP7Nepkqwpud/HfGpi9ZCi7pHonzI1KemdrRQU5CzVw1n+3R6a0q8WMkxJAc30L
WphJ+OlUwcTXnA9Ea7eYSFUCya52mihnYvBXiC91oLxdX/1q3EJBX26tJSesXUMs
j1ZQ1HJdWPNzFRteyj8xbZBhSWBXx+Qwx9ABptam1047xAETwFeMkWa2XsVX2cpt
OyC6iCNugBJaI6Fb6MQOQQ1/f5XdtdFsl2b8snhyYcwWj7UhFtbGfk0SZACtgrju
oVwwzmlMdvjK08dqQ29w9ybRVX5fRTrogw+jQqOa/I0N1t12yGduvESrzexRx1Gy
ADLeXPtqpsaU86di5mZl6nXZDqEQ3uZpyHEAA1UAHUiWV+QougYd35k2IpqENhM9
cokE2sDKPhi+R+sFweo8R8s40oUrjJtjEcP0wLngwjk6Ps6CraOx5TrFjkeDeaLL
bz3StAKxSs81HUWWRWa7eaH3Nl2Wu2yJBXOWfPDRP3lxxZvZfuZWP0peZhxqksBW
9mXldB7lbfRaAB50gy2G4gLKAAATugeFIszmSOJSwIUulbIczrYFd4m3xzfvz3TT
D/5avoCijczmZpRUprwf094WVA2Hm54TnT/wAIHvDeYPFPBHNFVds4FqTmyqNs6H
f8u1wfukMkAJUmL+OeXEsRwvrmEm4B3PAgJOJhr2e7oRycx74ULBegmupPGDBZZg
kpckSlVCBEikjlknUKXJvaubaiu5z9xn1gx0JkbsL90dWjrQfmZEY3YVgl7vvls9
yGm0QEEtMZX44+NokBbpI5whMbqW+y7IW74fzguWs/m8vqy1kexc5YfR1CiJgGYK
I3HtVTgjQm3MYktDEvFPtCVfSjbLt0EsFV27HGwkrioJjpXhIEB8SzCfWgsnHjY6
QUoJTQEdvbcoaT0UhJdxkBUqkhvgApX4k5KgvxIPgiKit5tGgeBwfinY0AmGkziS
28KPOaTgTBfgABNgKGfNbP4VaC+Ai/7BZnTCwGCFbeD3Tss50DrAhjfBoXMf7GcZ
T/sS+ix0kG5/xGhmmnOqr0tLxuhB9p1Q4GSlQd13NBG9kXfuJyo8GTMNGxkBHz0U
H2GjyiJ6F2UjoSGSTPPlRq9qGlBpWhdSGBgSUQLeykbLNgiUBCtjPkPwekM03rKq
PVEGARF3IYouUUf+naQzfKJagcfYByiv4sEkyOdKraNJbUZMl2XljEMRW52NSf2y
Q/c1JM2GqRs7YiGbUIdeAqJRHdkZOQbPYnX3LouZI9hm+M+nEfSKosUbeyGxpnXg
rU/CglxFJUSNi0fXXilDGpcSptphXtFSJAJm2f6J7JzHY9laXYKfaJLb/QxbFISP
kNX9X2iJ6BoeHRpvanmi8q+OA7PKjNS4oMBC2RjmPJPYhSINwEsRvSruczyYrcUB
QOGRwi0csX/mTzGmsKIr5+dybI1FPzciYutMWh418qQ3+tvfRAKXvUm82ImlMXbK
sw3Ix2rygvLgUBbc3/dtLhTgYtS0sY7Hayu0vqsdGcy6XscLNkoJiCInKV1+EDkf
wk5v1kWaSFrq1mY84pFHObrih3WW/eD5N4ObU1CtaknB3j0d+9WKP4o3cHJgwb51
He0KLDIaK+GvC/E8AEgR3g+gC5Tgs9u7WU6kWguS/vbDZ8JWOoUDJlgyRTEMp8oB
1vmxSpSo5kDzR+RTQIgiSzXVmThRVQY0vTH0106j4YotWb0BbBN9wMB97tSRo5t7
GfMkxW7Rk5rn+h5XutdlvcCjyyqePQ64zQtYamMTZ0InJoF9X4cOznzbvupCaEU3
BAUS1Lr30L7lwXE9WkcFWZKGQRoBgDwDc6p1g+lgk61c/LP9idoL+vUcck5EBL8t
IaV0yvKpVvdc/72AjAkJXmmidhZ4mnTEIwJRZmLHXVxXUndUFF8UT2oOQNuJNxim
M1jtgqGpIWjdxZid2Ap00cLrJZyH/GNYwZRxNnELfE5blD6JSzMrvFDcVyAD7r8n
RktYayXhm3Wr1sQGPe4lxXdTrcGGV10iLaO6PtsLWtc=
`pragma protect end_protected
