// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:52 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V4YtfRERRsQ+KyL1yRhl1U2GB06rAYEbJnxUAuaZJaTC9TspOXlzxCjLgXNrIP1b
KyG0BQHXZ0j83MDEYhRNDCjDldb71Fu2Jfvx+lLn4cxIpkRCw9h9QWpTbzSjAONy
n0n4tH9wTsejVqRYPg522Zo7f9bcWnIepubcE9q0b/I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30624)
JEtaMn61mn4WaRrDSfziAsoUl9ZO9C3ZQW2CVgm39XMn6G762O3QY2jM0QaGPiZV
fvSQ5ZpGA87cNvzTjWwc412yXFByH17mlsMnc4WWrNkrQffc1J54KhsmwNGSwQC6
Sv/v0PjwvkXh4evdx0VrGyNbAemvDX9AJ5VY8ew0c6DeKYJWR/CRHMB2ArlY4e3q
hHCOSUBGVhtVgq9z/Cu7XKzJSFihpzBIlvmQQFVK5wQW5MvtncqPt1BLrUgwUMnz
kko4BbZKWyZACV8ljWXLcZ5IS9RUz+jh40l5qVa77qR0145b1qIaZ+WgmAXG/XST
DGpntFSnHhDH36mnnn0w/NZnFrjygDVhN4P9Kj8Z89+dgRNwIrqPCJ8m13vMWyRn
RtgjemHmKAr/fagJbTYngwHp8WJf1xaRXhijwKTqYsnvxfCz84dOxsFrB3estSNw
IR0yNVsUamkdc1YtjRlmA0eTqzgSkteDu8gcadUP9Cg0y0C2h4oG+7gE1r0lTAtr
b8rxA09rW2ri318mbJJfmbfyiTqGAy46HcW2BQgYICp5dZrriwxXEsILCa/aNVWi
pNgYNHabBYZc+HTeLEhRc8yRhVPMt/3QGtC9LOWkSmLraPMMYxAwcXZruns1Lfnf
QJZPXypFgLTmF1V6IekLRx6Y2dFTVDbTEMhdz5yQm6a7uL6lW8xIqUTB/iYfRRQV
ZJfFZUcKUh1jKwA5YlsDvQ/Mgl82k+UTPTeoSPamlkGQ/HkslMf5t1sfEyXxaUTh
Lj43WlF5/nyHbtP0wAa3eMWpZ4tgwm6PImWOOJ0pMdSmI6NLIQ8l9q4S3zLQXFzf
gsNeF0Or1ZJD59i5J50qZvk6BnjRq2OYP7DkUZYtHSy6xCpDrG/aUnt7Rqss0dzh
f69e8T/su4oKZAuId0+17YZDN1zzd5j47HmGg0RnVMLI7TmU4YA3IcFpyhqC43Ev
+U1Uqh9/kCL08jxcL02w3mhoHOk7KFzCUbPFZJM6imtNHEOwLFDdmIE7V8wICZqZ
Q5vZbugzHPCnvJ2WPDoVUCyRVgnlnpP6SN+0FwqzGIzUv2aXrj5C4jqeIZx0W3lf
FnoDq81RQI1PKTBGcOFuTpUu8qa9FgmfJs+ZclG9MIWxanS6vNIv/V9p/Y5TLbWu
H7TEJs8g+hwWrnKYcUGBBXioizb554o5s1J0Txh2gKhGG380cjpCLCjtCN8/Ah5E
kk0cS4HNWW9KzzCObOkc+TPEu8pur/IysxMRiJ9L9RvAfmVv7lJFQ29y/ozFpmEu
mMSNoJ6bvkHBDcfG0YBn+s91DnjUHIkWgwu5Mj0h44YcS/peGFu7e9aINQL5vrph
m8qKSJvQ6bWrLvoHIJoumrKEPrqh9VBzVgSYsLGJht1WSNuMoDnYfgoSwTOvfod2
qJVkCXQdF4IPnqDtdM6lPjo1pOL8BMxbuqmhUPad+TkT2gO0vSuzV8/SYmAS6ttc
Q0P8r/w0ReF3qs4TzsrDrjQV2Aj+VFt19jkeKNgqTI3wO93ojkoWXkkDrap6mcap
lKvCu6sInrV75q7H8eCPbE+OxVZEtxsy92xOjecPZFe7Q6FpocubrH52KvrWX2Dq
8yVllLLGrRBXM42OR7wMXxi66tFVQ4hhdxCzEJXaxAIRVxyw3u9o829retxjTTbr
6S/XByRziS3u/5aMLCSJMyF+tAQhQ+Vi8nbJT14hAiHvrRGIhE/qHS5TQZmz1loY
AEaZDNhler8/qKXno/uQqUwDSmy+Fb03dByFIkxSLUoI5hB28txoihNGWxxRtM68
zN4uKcrDGoqWc44on5i7rJhUe2jy6nBX7UFUc3Bs4ad6pzwu6tAZgbFIztFwt5NZ
S+jRonEEYSBrntoNDmr/8cwqKUNjCp4FK9DQmyScJiFXqTGwef0aysBFffgenFBl
GT8f6wkEh+oHD/Zo+SAv0GfaArvDgy/o5T5kDBtZzU+XR9eRaIdtcjYCFQYw68X7
y8Ay2BpxjLTKEE1P4x22eVWwCaGdR44ibNebWFntB0a2FGobkYFiIg604k5aVGYK
Fef+Bn8Usf8+ph2UkijKZngFkwlrpN7q8ucxHYkGr+Panb6w5e7d0I21S56CTea7
F7sWxXTpFKbwQBkBG3uvVQmjy2gzT2drnCVt3FTKiQMPqaX9gfeC44nIZI4VugVq
BM5XAbqh93+/exgKPu664hxH4mqaAZZuV2Vg7+r4cfRbm6zTdvzFdmM8PalMmaGr
vsR8nOVOk6GNJGokT+mu0RIWI9a50B4bE3TnF2m46G8NdToBvK9MvEMCKvxgBovQ
ZZr+JQEkDgd9dhDnuatrl0Y75JBToD5pdbfOAxadK1spy9R1jJulJoBO5KB35yVh
NtXSbNVT/Y8fxgNBRaJpj6yEod1NSSss4Ts+EWRFEpOZb8tPRmi7Ocq9WHFuGvWQ
z8A5dArArcklyqeNVWU1rt8MkW2EnbNFPAch11/a5SbV3GFDZD9A5A3de/99lueP
ZQsTgfUz5DIxPLmQ0QzcsSj3U4FAtrDb2TFpT/tp7zFoeA7X1j433O0lU9LKYVah
ejZAxRDi0bNODLl3+Bw4X3NIlSGXXNyAICXHsvzbNmjzTJQZCGb08gitUIDAPeCi
OLa1m81jCzmGnuF/eWf+6+JcJHzhY7QO8RF8V1SrCF40zAj817LWItpxCjL1z+LP
0ccx6GcXKCm9MfbmfgBuL4Uh3NaZ2EMK9iyKIqNTm5x3eoiVgijDV9LbNd9pY6Qi
XElwECH84X8OAnBsn+Ex+WFY9O8qVwQrT7O9pg39MIYKkpz1iD2gcg77QwQZS0lF
De8vZU4HE8iYCkk/8FQ5yTbjVuMX+QG1UEv+Doy22IIhYvHZv3wS+67lpyjzTfkl
uVY6btYDLlN2oiVAF2xTBD/WUjC7nmxk+N71qKY2u+N5zBf1Nz+dJWmPK4cNYXvX
3m1+lWZ1JtIpg2OwrBEL8GWBU4olCCT8JRYKAJJrC8maMFaBR2fG2lhxW4suYpu+
AK2aI23NtLY2gWnWeT9++hycQW4/Yp9Vy7H6LOBuQqlZGa5YCQIUrlJVlfzDKv6C
eQlNJzto+aiN0hy3YLHYdWO5txnpECYL6D93nWH+gkiq+NpOmUm6/mEb9V1Fwpai
ir2fN1t72wccG3Be+hf4bwr0RmEQdhBtRIONMy2KCOj/S5DIWc7AtdLIzmvYtkJs
Hnft1+pkGWcL5dIKEvlPph3NjQK2wve3LtLXZZ5YRcM3OWjhcq+HDgHF85wHOB7v
sifvj/c7wdME7xFpfxpQyH/v1e23HeLmWr8jkhpWewXpz1YwVJTFebZhyYXlyf+y
WSrOcrI/wFUXtgE1TIYxKYCf5BWABP1OIe8MFuOsjvY4PWjKnFnOzWpCuPmAGUi7
oj2t7ISsAFbDMkljCh045+KQ3JRfTp80xvVP/Q123Hwa8zoZkhOYdvJ3xCmfbjqM
/7tN9GZ/DzOO7gy3nvgFvjGyufy50bgAvmfoTb20t2vbSgVUbwipn3CTNICwXC1i
VnMHtoiJsFZRFdqPE18oAo0C0ImhZzUzgVQd3bZrRoDIJEXFTcIP7v5NEP4IeZ9C
DySU8/n93ANWmE/SD6SunxbPAHKZJWLXcZ+EKTfSkvU9GDcM4jynKXrqvxODTEhh
2YJKwdA+QwixBZVJ/I3dEQplREXFRlIJs0rG3vNOS21PrVVi/oUDfJPjm1mzbk9R
WfoPa3oAiqBq3IRatbsiBzLZQATzPQ4H36JoqmjbA3vPagunn9oD+BVwmNQ41gpT
13Iyz2XtZBrTWrU8ZnFB6bNTz0EPtQRpMipbK8hPaVbRfY6k1TqYj7NDO1d7sDiD
ElweTOcYbIfYFweud7RszLRohQy4dg7mFfSJiMExHToVT/euOTck4zC3Jh/v5wkb
/Dp1SnzgfJoNQdwnnGgDqOzFmQTTfPWJqXisOJFs9ztE7ahsCoXI2QxSbNnKG9FK
9xtdbz0ytvdnRkLGfRdbP/o1BySQUoBawu1xricgb3Gtmu4d3lNprOscL2VVOsAm
9Rl/26l6GX58NkcmT2pItbHYRLiu5OhWD6II+KhkREO4dqazg5qtKlFvZySGxbxF
073aZ234TvjijMp02hTNYhB5hmyUhUU+GK/FOMb9KnyT94Ef2WE1wzH63bbSoqcn
AORlfVaXvs35F3bcCiu2wyYUeWBruQraU9vdOJ95tH1w1KgmbNmU3BzSft2qRvcR
p86DK3lSAbl4VCS8TLQ9UsKS7cxyU/AqzYTx1Gu79nTE+J33ogMGI9NnJA4WLPY0
NzonzkbSW6F4bPIJuo5JQKOFRQgt4HUCMz0GNRDglcJZZczeso4+z26coGWg2vPc
w2yr/rQEAyaBI45erMEZlJnLxmvWRGFFnngP67BZTw+sftdIPNS9w5og41Vy24Fj
IxdvhTDs+BLMvG+Dewc4gT5TjbD8tsAWKdcmS2yIfTp7uSPMxhY+lFtCOgAvA6+g
xeUZnqffhrQW2J8zIX2OWL574ZpPgHJBNgoJ9cquQuLXMOsRYON5zt66tbGrNMiL
/PmMDLNmE3i8w8jqtHkiULCQdOisYySeehoQrLUlINvC+hOR2KBkpDw8FJ29i2Rx
P6aemrAYbvJb5wh7G6tsUrYhjphAyR2Zyxt1PrK41c6BGtDXeVCKc+6ssNgfhxnQ
AZG+y7E9OayjhwP7z+n3yscCAA+Jg2uOgXxjh3LHiqdSFPqDCuxlDCcbytMgu6qO
rPDy8BYJ6K+80aSEMFG8DcoASbiA4vVllz8DJCRz3UiNnknLeYSLw68iN/N7SW4j
I047pu+uvK1S7vaUZFYPgYfs5wUVHPD/pi/BSQBJThOalt90dxYdw52cJQeJA23J
hU+RASUkRXnfNCLajxPjwUxZL9x18X6LIJVk/a5HaKWaJi25ddFvEHZY4/IOnxD1
obhAN4w2QRm3R1Mknti3GalI+Kv+2FC5ZJKFQZ8fIMf1fRhOeLxZDD4YTRZGRUDk
jSySHKeMYTu85IEosaiJxrEuOwTBUGzdVkhUYfjy30ExkHpblWMilfzIseHboJ4E
u4RCrRNXRvcYF4BJoilaD0WtkGMHgdbK44Sxd41gnv40qY7lXjovDBNsPBv/dY8l
KqpLNZRcvmeC7q9gVbZdo04jw9QNAc5c2hMu1VWyqd4nPwbcDihFfwH/1PCB7Z2H
JGn7qNkBcv2lJXpniXSM3EP83/9PU5RrG2SqVmKKBQE3h/MwcQBiG+e9D3EfHFFc
5HG2ZxFSCh8DIJ8L8rtQfAgt+70L3OsRnSmAJ54Hvh7k2aO2/Z7Ww27nQOD6DCje
0xivzuJxsGzmMl3YzeQ4cuq5XGvFDCuVK/ECIZX0ZrZmOxOamT2qyhg91Clk+1Cn
aM54XEcjDkjG1FJFXg1dqVrOnQ5IieyxFGeHzlsOFXkY4S4b7cFV4qUOrhroBhSx
kDIzcMpVQrkPSMo/sXRHsGXtTevuFPd8q8cscSqTrxkI955hnCUgidXr1O6OJVnc
lxH/tS+HWm3pmB0si7krZXdwr42VWTdicJEnYd2dtEl1v4DpjBQRmijRQm6uKD1B
rezFb46nLM6M93HBQ+kov9j8Cfm9wygegsoTDp5Mu/BzOW+Ub2nlTSdP4L5jWZVh
4lGLBeh6p45eaDsjGieKD4wcxi9Ezd+R4fArGUhNsIJtx1XsCKZXZKF/j2RGoMps
TZos6iDMwINnZXk+MrWOI5N4Zdj10ivkX5QMv7f96SOB6/hMl4h61husQloxEunC
SdHSbc9wtuxcj63b3OYbYfhjj5Yc3UiDu5Tg4dI2IPjsYAGjLmHILeHVxjJ+MPSE
i/PyKUp4QUFTX4rfQ/8faxtfStDa2DDCHH4WRebA8K4CE50lsCAFip0NRawkpWAX
qawL2JYqo77ZeRsmAFRV0ndC/NDuL3bO77826AQaww+VVRxmR6ph4/SdzRoWnhs0
4D0SeOleIGJd6IDBQqH/1K7c3nqso6L56Wj0ZevJBw0lwtte22hHkGmN0V62UQS0
lGcfWx73yhVDBoE9NsdhUqRqKcRk6qPfh3dw6gWvm4qEB+/U0w83KawZ2kFsnnr4
4mm3HsX2JeUS7UXrm9YsokidhrUtgKX/AX3jNJGwI0vzY5fQKfj3OxwQhTY2nO+a
QHMmcmJZ9K0XYJc9BXd2vNss1RtvaEXgvAMwQPvWitMY7q6PGkTx8xrDaJwCXSFK
7mVzN3xI17jcdi9DyoEFOU6siR8qYbVXUdQ92SkF/ocdtwwIMzUt9FtKEbhEebbw
pAwDjvvUvuQVyMf2ZS7LpOud4gj22Byjfc53eUU5PYJ5YdWXvRxE2T2SFq54ncSc
hSLc4cFyvVOkbfl2oISfz9XK/c6yBx1MYjEWyIfWegTP0Z0331FZ4jm4ac+Xkatp
7ACBA2m1yFQ2fKrocEadFriX6n7ND5tpe9CecU6PUEx1+tHWK2hCk2O/DoetOYJk
qqz3itFBXP4gUxDjXC1gdHCh6MQm+zY0Gum/+/CCqZ8uYpHJtXoaA97/rkjYq8jW
JhWQeBHf642s9gXnk/ViqImQlRcK0gWsCPQZVMGTBZ/WBmjMTF7cc3W4BHtQT9O+
ACOgLeW1jcWsWvaLMHuZaZjvweGFlrm9qhfVn7dRGRwN1wtZVKmPBukjrcCk3Kzd
+L3WgrugCSscAEBSx6pQQLot6kIh1dOSki+TSfcIKs6ROttFwUfr3X78xCaxcQ30
OA/Zeq3QkBrVBYMbfIzaF1TjhSUp/Sa4xfr+DwstsZpRsGzfg6dsNG94M9RpJ+ea
0J2WiFYWKsd3ymDmJJWQAXB3ZbG8agOJZ5goCDFueN1TbwxSXczCr3J/trtpgKfU
nmg4pdyU4UWRWVYCJBlkKsTBvyVCE4q4X5ijqXfONsAIc0++4gMccj6DHsyAfcpk
Qi5J1wyWszRW3V7MI+45aswrUmPo/0n+iqcyznNAuYPPXD1Zh6LjagY5tljoOBnz
hUNiQoK7ERwScpS0zqqXldf/rXVgum/CPXxl+I/S3iRQcnhzMjkzMbc6+tQALNOy
XFDBJMav+Ldx+sPqFakqSXScqOgzEmoqCOwQ8iYTPOZjvpqMhIsGOM+Jq69WGLK9
8nwFudy625x7WX6IBK3g7Yo66cH9tTJPYyHKGLKZuCBfEVb/l0WQxpDGtbFewebS
QzVrdmz1gXlVObTXDcAnEkX8mIzQZqqbKRPIQroRbOROAv+kYbtZcri+XS+iewgv
w0jf3RzSfRCZAm3U9Dmt3JHLfcHyj6TJjK66nhpV41J3rD7LsG4C1SpvIkH6iqfj
Kk2fVHv6WhZsIWI55ykvBmk2GYxxxTY0vYJRV+iW+qj9bkh2+gg5fAQP1j3NjB7g
Guz+ShZrcMeaLMnmKgNf7rFEdifiM7jQZlkN9Xp2g3uFbu71DHMrPmpJ574Zxz9w
/v63opUEmb2R1uYd1ilQMUk7HiQGorpPs5v0lJalVr6Hvb26N+JD3Np4dRLBSfL/
hjq5MnqQkzh2Rw6GC82yryeVIkD/Ab+V6wxw7y71OFES8VYliCq8ogUf2fvg49UZ
oB/xhd3VTv08taEfJJTpFK2/4RFQp3bKsVd5KcdAyHkvXduoXabqUxWwq10Glzty
dKW7nb3mVJL8ucXcTuimpqU9OzkmVpS7B6x9KzITRfLYuWW1fecrPHySC+HU/8Gu
fgGCPHSoYfKWwq13RtwJ8fARFubJhmeJnAIuybuO95mYiR1URStpBiHouS77NTco
vs6KzTO82Hj2VsWiEubrKmzgTzd409X5oK9sRCdMjv+CsbTt4euodhkE2nWGj3mt
3lFMIYj/XpHIx/BGjdZMdHVnHM1X1HdhBUm4HlR2uSnM1Ix7YDkTmRwI3rhES9cz
aNUDKvNz0thRAuLR1GJlC1Xz8FF47Wy6KiZQZHrV63AgDdchxka69WpxvhpSRbPG
vXR3ZwWsl6FC7PN423/ztmnac2x9VewDb6hNCzfddB9exMpc0EjZKpmMLg3HL/ng
FFvvyF6UpHn552TugwnXJa3znhadia8DPU7LszpyAWJXP9gEA9bPZpJoG5ZweYxG
t047+KHT4MgeIj9h3dP19KwjnGAZIwc0AGOtaodnI3vcVlsy8r/iMD/hAfmYg3nD
kbYlABrbX3p8Q07ikDOtbAg6wYPHNzulppyOzonSln69iMnK90hQ5PNclJ0gAbGY
ANZ5F325O7EsE58uBuk1O9QAZIcEojHitXJFpfxV4G6/3hKC92e1RS7FxRu0Fe+t
mUNO2840jYYuE1jUlpq9bNmQ2q/YHjOW/b5tR3ARLQTU9ETfJJdNXkMXLGMCzZgv
DMQQuI2ZXsizeew083btgCIdO/ZSXleCg+zVXjGk6pnJ62jSB/59vJrC5hC4qIng
ONhoakxpHBeKex0qh2SOO3jQCMVXSRHkrJHgA6ns5wqS7BHL1BNSQuBCujKIRdK6
Kmv459EeofkOBubQ+u0AZajW70n1/HM5515og2Clb14v377wtYe0jvRLGNxQoTSv
HKpEwCmCqPImn8WGu7KFr327rWIzYlPWEwqz5zn3jBWPPgnNywnafSI7q6g4yeey
c0LWigHdvTc0ZxbcguaZ7nE+HmjdPkKbUSc24Pp5MrIVBPR2IikL0GPwfOxQhSxm
Q6e2rvX3iKa2k0WR5g58keg0yJdAosOZj8uyVnZMpXw03lasFyBhawS+x+6lE3yJ
pfM+kpOKE8yrfbwgx7DPB6mCsekGmnukg6C8c05c6j3n9wItyYSa2MDwxI7iJ+jE
LjdUpRK9zsQqil7Rw2sqLlebwfgPTkQt4+1dfFzUUyLyP1jAg6UC4M0nHWmiR2fc
lv0iIpouLfw86JI9r1MItbEUyirfXsBAC/UvZDmXCVdzC2i4zNTQvN+dDI/U71hS
05BXaMLLVze1w64BPXtscLJUOQpUKIyQFwYJDes40HkwZeZrkwy465hr++O8gc8k
a2/pf77gZooI4kw0UEE42QAIK4yAiNEm8gmT9P9GPyWWbxpv5lQaz+r02255SZBR
WsSWOuRRrKhzAZz9qPztm1Rwu0ta2JMc195GeW7eWFSnomjjz49e77Sgy9LMTDsh
Gb6iYqki/mpq+vqZ4/NgjKFL5mlFtrAMpnhe7aWTopXyNnYbQhKTzOp5AiorE/B7
a1bhE2ZnjnG59yvhttc9M5+UCpKl3l4g3PhMgoicArLTkGZsTbttDDG5m8ptXKPW
vhhAMVIqyvBMPCW1Ki3R1OBaO8dr+MIscr1R4zDAJLmQya1bUwgW/PNf7ko3FOLt
ETRdtH+G5OvrA/zbj8AikjrZwWLewUC9LPoVpw6wb0eTE7u9lhx87F0Gi0tIt+Gn
E2eJa4PDaEH7DOniMDYqp/Aev3xa5314xnqiCsPtjl2mGxVZ23WeqtkJZ+JT/6i5
x18+PZVpoUFMmmKFbhO+6ixC23IK58fBxc+SOC7YJZvZzChML7tbMA/MigmwI0ef
38TZwlx0avK4P/tSYcSfGbIj1mpJV1bVGHwjCGtYfkEPGCHDysJKeaKDtow20FSg
4Sl/m6vU/5lsYayTnp8T9462KUssm6V6lhQ2v//GX/xEqrIr+DPdHxKUekhk4SC6
FdiBrbWU47LyAQHJFGp9p/dU4qOY16pyZKl0HOjagEkmlTHOJYx0HOpYVC/ZORB8
MzWwDHYxWdy5TMa+Mt3SMeACr1cOgbkR/Lglqn+A97FJ28Gw4JZMWW1tRbdAL77D
o2NBadyjU/Y46SQwgZqGgRriCgG/mHqX9aasWHTHU+RMkozWql7hNcl5YhsWi9tr
QgbgMKqfky0ccP5PiLodzeF3DRRQdcwPDQhUnhHNKx7N8TfHyCjUoImvh6Uk4JwQ
UJhcTsBOqmW/V134TAPHrbuAZltz86jwgr0s4okBBjF2JRHi/r5/E3paUXpptuy3
m3dwmzA/FSGMsUOaYo5GZXME3kcqP0NowkA4qJdQflTKD6qb/Q+I4XEcLTMseN58
sBNuz4GaPXop+Qqfe6sKimb/cjE2gJ1089zwDz/9M3xBzHLeAuq+TEHGzKjAb8QJ
vo3vijkHjhozhgTjA4SNX3QVB/Bdhnu5YLlS/WNfNBJmbeWKv2IvqeHGkh/UNRZT
Cpf4vZY10iW0/SWxk0F/eoSLhHFc9Bjqr8ca/B3QktHFQl+QPYjJRf1i+THX1wiY
5kwswLZgXyqpf1YoO+9ZlAVwHWXMNoaIVBlWR7RV0swIVDdWldbY9aOBuK+4+Wj8
fREQJLCcQvzv9afbZvZ76bma2CKuYAf8oK3LS5KN8hDDUCyfTgC+beXd0Bvng9D/
dyDWaM2PiiwbME8ornhAh3NVu7m30Iw22qCzXqmmVwwyScp5smiFwOl79g9rVOEl
BWukAZvwy38I+ZnX/RPlai7rRV2sck0QJRBX/FZfhLnJUh43fbmULJGtFZSXm5Qi
4CnE2RhayRPEn0xIpQd2+3DljLIQtk2hre5dX4KpoqnPfq0jyM2Vgcemc/4PyoUu
6EcwaWOqGFUl7m7OqMvUv0h9nu5DZMi5YlVyXb3+yK61YNeD8/INcT/jSKBqA/vv
hnSxS4NBhfG7k15dKd6pXjZFvNBJ2FFAH0EzgouEhDU2OBxK/fZWnT5iIphGzDH4
YnvZcT1aY3ZLme2WcAzrf5lk57UluveNos9AgMgqEPQ1tTta1Ax3b+WtvfvRhjMb
OqcTi7KeI0hG6SX4JDS3oEjKFpfoqhvsbZBwsHZG8P5PSxavfc1gUCAFIKpApxQL
lUi/3/dZi/2b14n1AoUsZs80AgUZVmxiRAMuiw7Jeq3ULN8bH/02UKlDv1jxKlso
/nfsWzWh4sRHQFGxUZvNsZiXKCc7Tkj+30QZt7T/NHvYrFCBB/EytbKuGh9QkAy3
Rnn3uRxsdsfYT4LxBFk55VX+Uc5n9+J38o2U7CT9abGhpaQAAXSkL2rh2mdr613N
dtujbLZIYLshP4CxgPhMI9KFSvlpfIM44Z00Db9cxQjxLtigJTyPc4MzD5Wo4nWL
0zZ6COPNVtFTK0g9aQ08+E8/DJ2gfS8zpUMLRs9dTf5s8pVL5cXkHeWSFxUR6eTb
vRJ2bruDLCKetA3bqMeiwEfEqZVLoydwb/jRs8E4Jx5CmKNd21x8v0jkkif4LCgG
ZnTsNbDn4RJl8mJAzNugTqmkPs5irvS9oXmptPI7wvgRlode7w/xwYM0wLlRtRin
cbi9aaQ7R68cLtuR0U+gNNlHiGIguHiGGc2ZnSKJl/u32llQpFgBbjimG1Ws8Y3K
wvAnt1BceeSyDK1DBgW1PNVaussWqxy18VY2y70TCzpjlznvtDNPPGsNYhRA7ih1
pgwmYG1y0K7QfQQDpoxzU9YSDklcXCK5QiHA6vYxPSEzMP71un/hc8OXbjpmQEgk
eT88YhnrAdhkqncX2wbT2ts/K99VnjRu02OFTtl3y7yDppbDfcnq1/pyJdZAMESm
LSdnsA8zAE5jfAQ//1A7AMMqv4E5AJeaOiSqg/s28FpNuWKcvbd/gxa8BUHlapIu
HVRK1TuCnj2f8wVIjHFUq11dz/wLinY1rMZ7fATFBNRRu/Etvx+M0hcnl7BLQEpU
tcYT3jH7J4M/8/r6vhS5tWSECxYw1eK1UBtnLTT/ITlr5tVD/glggiGhbkJHb5YK
4rpIJgGDORAOpmcix5wiDQqNepPZ7B3XtmhhxAqF7BSUZapoqS2FIYWdusvzC4bh
BOvw0cP8LzEGcFKpvFOvfPZJc/84DnMD3mS9fcIZJhhvUk1C0ho9UmniIv+Aj4VL
lOtpRtG6bMadyRKg/RrmsDWkM+Jp/esOY+d50+65StKvQMJfZwjfiYz3RB+NdMHV
sFiO9D+5TyIpMp2HEJNZ0qeAY5uc2l20xfFhKpwVQ4UL1J3M7qmFYQ4jRRX6kF9E
dA2xZhVKIdZ1lRx6OpXa3T7XV8u0u4rIhKioCluZxcz0cRfv/gHGmS3cO+NNLq8X
tmcCg3juCe1xJqCYThCwdIs1hUROjX/iZCrwJNyxPm389nS7c4FxlcAL0OPRh1dW
MQ5Ud1MppKj+CykM3Og3mZZ+HtFcL8aj6owLflOuK9aUdqm/mqcf5KMLYPbCmnc6
pPLh7G9WKp9z+oiHmXdDcTMPNW2JcT7kCKLisQUM9SdLNedlOOCEdRmdL80Vyek4
+gClf3DRohnWs8p2gxhJXWxQZjUw6VZVFyz9wm2xq3z7vBkDiL248WD+m6o2YRpc
NofwgEUvgsS2QpD41l260lIdHmr8DT0NoCDHDlAFqkfE8eA+KJed4q33g4eS4nCj
Ev5hRRi6E+0dtlGLyvU7X2NQgmKYwMe+ZeF+4V4O51nh0cggIIkF9nFzx/vuGepL
Ex3lSyIIxDqdhoAzZFB8NwiTeKM6H1A8a0rMmywFKkxzU/nep1NTLX20st/qx6AM
9Y1W+VF4TwZlC9qIDsfFMEfyTKYy7u36R6gVewtDSRCN3qAq0DHyIgmEbzYc09UL
4m/EjF0vv/IkBriqRv2fhv54t8AKJHTWQ6ZoHgUZH+hgcr2b7+ALQkJOUzijHxkj
o3OJNoN08GmKeb7uU3ugrSWE6wZmrQfnXIzVUXyCGl9ty80gmtQZk/iiNhZYU+cW
KNwKVkBynmkIes5oEQQE9oGcwepQwiGvaHThaauVguRAiPQR3A23118O7PwmM/+c
SkYsUTLk/iU25WRny8lUK4GZ6HqSOqBXyIzdFkv6UNzzZjhbrJ2jJoVjN04ZnXtQ
xFLIi3+1Hmtcix+GX5Tj8wgtWL4ieRFsqpQ4w2lboFDIS5o9q5qTvGro3j5zgnUd
Jllp6vBS5S8o0I7B3RyM1V5HA7lX8tD6rCMKfEd0jJhCExyed+/zWShNH7x6NTH9
queNZgo2L+kXjpWzDYq90Q/oS1tOf208Get92oibJ19HrxAf3w6iUYLB6+/bo4Eh
qiWTfgexrEgMBV08xQHrUJSH4fToijfS977UnzCv4LwEMNmUxE7ADYyx6pcB3CA1
R+izRM9IJIqC1oQ+Lfw3skbCfMj2gvtYxm9RZrMLBZrCA6nHc7IMuT/kTs4y7dhF
17/dYJGVeS5R2H2cfGn2k1BPdnPGNQv2yj64GVPrqsAiQxf3aUpKBLUzS+MfJbGN
LzhEEnqpp9k1IKcto29k/K6e4HHlfETJl4H3afCN7rHLb1BJCg/qQ7S45uQAiNgb
F8wNzYAVgjWiAwbKtLviop0nqNhzHT3Pt5k1TJFdYLmB7tOu+9nj8XtSAIUwQVyp
6nFP4DXZUv1sMiii88UTNW9DwGzt4JWChDkKlu/P5cHYgp+OrimRNXhDVjOCh9To
LNQ7cRBpTLd5T5c4rWXRwKPRIWMZT4N2S8aJ5QuDZtm99PxWiwdbqLyCzUo78NWT
xSpZD8u3QykmOSiqcbcym/D2UBEg2wD1m3CUp7h7zv7lezKqolpI+HN4S+BcGaY/
ULDwcm0+9EoXjinP/Nge2HPaGzM9TL2KvCrYVty+bWXTJVqzSgRv1/fUvu+8y+H6
YpIh113Q2m7GPnAaPj9chklq2kjdoYdo6tFcPisO7cg5kXgXZilqBDaB2ZfUynuj
Cz4wIMmNTx2y8bk7paeiDKtGCCXb44ox9ezejbfSFryN0MWddlgOXwgzseJT31n6
Jfdh8hobJMjDe19/0J1u1bSaqblWlyJUbdU6mXekpt58RnjHOLs1dOE6n1uxXI44
Bfg3lz2JX3rDtCL02UDbTFPeyvx6ZdMKfH26w8M2O0zjGDzHtdtCtPmi1qk7+LR7
k2yKGncAcX6bW6dkGCW2IKmT2WjcwXJcOkDvUjpzWs/XqN44m+hBWj/eNYucA0p2
0gduZtl3Erl10naBdkqOgCr2HAq2rqhQ1N/yMw+d/f5x7pDGjHThVZAqlbuRXcSE
8NL0nElN5pJITqMW6aauxbcWhdqszLXLBlMGbqAcJ7HG0cFIryt3mj88McIE8WZF
5iqfXqY5PkI4qOYMhlzvmuMD0E/UKyxi3Xc4hCddXZwfWcsiqpLmUHG+BhYSa71s
NK2D6Nyt7BGu7+jRlMO0sPqFKYUpKfS9BKncNNe+9BlzIpGijYj3zzRwlIOWMdwk
lV0E80KzUJTpA4HmTR1MgLrWTISrZNuYtCLjBjhdVIHBs7rW2sSKhMXf7zlYLVFl
qDPiDHhDOXCGniyF6D4rOrAvuHqxlsyB6Cq2dtY7VSyF98caictGYT7b1jejebP/
emVYEHGVm+FrAJVBm50mhEi5UY8SpnoB++nNzTjQ97i94+TeHLnACCVACtgEI1jF
HoR5Wmd7XcBV4AslEXGm9FTCl2xKOOW/4adsLl7eerhbRGJLLDIyeNKIH72yRBv6
Xjp0Z47MTT7dVsHBI/9QxmFw0UrXgQt38EDIt6Px6gqb1Q8pTthX6FjyV4pImAgW
e8LMFVOA6vVci16OaZGQT23lwohCt3jaQLP2bzu+Dye3GXNnkkB4fwzD8p5LAvmi
vGkQGgVuYZWaPVc7R30KbttQKm15MIs2o7GYJdQBmk5xeL5GZc7DsDgJeYzPQiE1
OLtwaHKxGBW1Kl1NHrDNPn+UozKPAGeuoHc1XFD/fu0Zc41NQdS4Z9ulADsMcs5Z
9Gr9c0J5cvQxlugbB6BVnV6Z5eLnOyLyriQSqlA86k9Vp4gfUFw7F8Gn/4NveQpx
sFnku4gtJQ3X4BsFPrfyUPD/MyRji3Q31vD5qNcJMpEOBqwO6ylf2Dwmjwg7DwEm
fCpmrJ1r3b3taOhrQuKRi8XxtiXvwHZ7fB2JF2kw5fL/FNLYDVB/qL3sLfw2L7xo
Wn3LCrPi7GwuSQuP6qqIbS+5JeMO7y/vUkl9vvIbyPoC+njJ+hytRySOU1tXPdHQ
hhDYaS9hta1MK+mZ+YtkDPi3x4A+NoU5nAWM3euH4AdHi8VCuMRrgFtge4zxg/Em
2WrN3kB4RiFYRXC/g4Lba5yNjIazkrqSwgBDtImt1m39MT3elcGMQcSTdS6WC6+l
0we+dSjVlBsZvFFh6STsQ6Jw8zqxAfjrZxT9xAEsXIkMe2wZ4+PXye4DMsnJxF0P
JHC1FMg115WQ7scTIW8L7g09g/SBWU+YUIGr+3sZZbbk2cnvbF5CZToTRyCcsDt5
Q6+wc/L9o+lBbYqtbVLOd9I70SqGGos9a/j04YylunKiVKNTTaYJhEd5cVDlBb/W
b3HNb25epAtsnrhji32Gm1t7/r17lMYjYFssSdkrafIHKWYrWMHHyrhUWrCaViYa
vz7wu1/AeOI4KBu1itNcv7IIrbHLj32zGQxdoZs93YwV4Z9FpC5EjDcdJ1beGl/M
2vFcMBdlckFY8MalwePYFad6m7zzNB9RNlfQi0FYdg0FL/K0CF+DzasDqay/zuL9
1fImnkDmhO3u1/zbeVbOiG9kDmbXTDzQVcD5nFr5o4Jg9l9vqXg1RQBFFnPr9lFd
d8UzUnGwsGrXlbxXTgY9Vy2c4xJX20wOPugAhdVgaSVkU+KCbSZbcQJRt3WAdMZk
jvZyeWyYs6/KmOKLNcaJG8hAOnJCnkgjPYNSj9S/ki0f4+4JMFo8w7rr6n0Yu2hE
4xf6m/KszG5/loNzZOohmeMQgbLdORapvqnzvfWxVizygeMfGzZe3fokiMsWLy8p
x/inJYin03af00HpxoRphUc2NgDLsUoWoDcUxN285a6FuoXRmUp0+Woq92R/voCd
k8gc8yacsG58kxbtPvAhOSPCfqfNrEl0h0THE9B6zaslqcBoOm76qChveF+XNr0Y
rQfbBJk3dLP1qFChRGnmXccced6znbLwatBseDa/PnmJFmWjlLisP2Fv99HpuI20
SEXVHUSJR7B87/jC9WM4vd6/WpyQR/iA48xtxlQ4W6e4u+vYPk+W841dKZQlqHxf
Y4zuCp3PH7jYhMakdqIZktlHudCDQqSs4cCITBGm0e1bHvA67PoJRsDIwKG9UvHN
47gqZFtIrZ0Yov6h2J3imB9wSHa2SqahOhUq09XLqc64ee77rTjSZMhdxSQ+YTih
Pz8gSR8zQtsIjeKh50g9gUPz+Q6UA7W1EuUzGgf0B9OPe/NU6icmJ1xjzmdcsL7y
Jm3ePQKhY+3vW6eELTFcrGqNxa3L4sZzM+9BrLvlQxfDQ8RecWGXNwLHmly4aQa4
UJI8VPUJ9u3vFa/6W7CCxsYPRfUnnhsX2dqqkrUBz2rR2aDnXlTO0NrecoYMpqMN
DRPS2KzvUzFEdVT7dVGfIUUAvPhtFwEaRKi4rKpZznkSqnGGJCChcJgdUZ9N8pqW
PiS7D2Xziz6ZYcftOy+UmJkINBNLYW/2NEA2HwKB2MzxhLmci57p699cHkIHaAZI
l+q+d4etgaq+YhxY0yInFwLGQWX2nc6O8BzkR6y6pqoOwyCSwPQNHl0eHveE1mPu
/Uj3PMtxS1+1Bcx0bl0zJPWJ6daqLDVRFQJvBEno+TJBYhb+zTsF2ULJ88Flixf8
irXISGUKli4TyB8ziXiAxdVFBZZfuRsgulk6GT0jT5IJ9VQOz/NLN4T0jce+PFqz
H7N/vFbleqh+BAp4piudi7Me1O1W1kv8swSzMaXeW8p11YI0zZF5ubyxE0isgTz7
oYOHwYMY+iv5Cb8eQAUFG/u56vrMrQlUhYCZ96I5Bc2h3AMp5maQB2WQxtxaYD1n
xK+0+oZwMDioNQ3IEMJsGqs1TEuKL6yPrJ5A7PFKObSkBRwetmfH3Q+ljLIRJLg6
J2mH0NXYtkzWl7dwmPCpxZx+kMZMuNGsfNZGkgwS4VMK7Vg2vD/fXDuPwrlQRfaE
N3ze3f+ukYYimIEagIjd9lKwxQK3Xb56qYF/cjGnW5IkKWgg7xXULqt6/dQQOUme
7IaEJFFSuKxX7848lXqbeg4dSp6DSXkwyyyg4eKcg+3CRq2ht+HRd675nIt6OAmM
ISXHxdWvl7xVkl6Gu4djf6WOFqNrmvkXbrrtfO5OSAVGQp+722Q96SP9kubunJwk
Rk0qTJuFmCE0Y/09SZLvvtT+sqIT2Y+wjyxw1O23wp9VrOVg8lITWIy51KF13oUG
gmhFMM2We7+yn4Uibhhs9KhKH1GEUzF7S6ZHQkukTuWltJwSya3cuL0Ldzg1+bjp
dx8XgIHB0be1EqYesr/NJzxzY6mvlVB9x4jT7xoSv/4Il4H3+B4QmAwgKgbP2tfp
FDJVg9WvZALxpWFmFwQ7GpdFj9PZ6juk8Ho9mpfzTfrd94pvA/x+e/70HePC+8hY
8rFMURU8kEWTyvZmJulxvHPqhSrnA5SxBjLSzLqG/fYlL1/HXL4a3wWJ0lOoIeLr
VLN/YFALQ5k9JvcNeiHhroJLGc3qX2V6dUI/MiS6B1m+XDRMrxW8LG0cBP1ifUVz
ZMN2L2X/2WG250V7unC/Cb2vGRpiLMllNUJddbbW/8gFT52IvvGcdV5kIq6bANWw
RBlkqNr5IPlYPDVCXMTG9NozT2+E1DTPk7RfBpZOUshNnSa23jVzW7HmJX14t/sw
sBtqlSF0+SBH0+5iLSnNnfCXSE0u/e2++arx4Qh1m4T/1GqD3+7xl4tiKF++ApS+
LuHnNWEgHIxVfIhXg4iHZEaMSwHecmNbL3f8bJoR4MHLAFaEMDLOyTy8H06v5G1z
0e2LCVruMPCl83PxFsraxO8uETIjId05hnTsDgUAIDOBqzeDhiP4tjnY/J8aGiff
AWrIuQSYeTjBJC54Ojy6RwhmsB3OcIVENmioB4KNmG0POjii+wBq1IRO1dwz5O6O
Yle0ff8l5cy/Ze7eZtruJ1eMSNLRejL9+0RX/qQVDscz74Iizbg/i2lciW+glC89
cyt8N9JmVbDIY4qSMMBBhcpVaKwskivfwxTrN42V4WhwAQ8hcoCT2nz7j7gbqdXR
wBb858T098N8UXsV7bCpBLuvlk1y/v8WvHIUxujPa6i5BRzD8+yfOpzOZYS772og
VQqO7D+ZBjJ9TaAQ4a2bj5UwpI6lsau05LcXK/loHqffatQByldPh1hdxTNABU2R
/L8SFk4dv3a+5mjEWIUwKolXOI1RAVRmdqaw9q9hOjq+yoE5B7wPCfB5HhWW1JDt
40eJRDSZpOj/op8jNgD45RVnhC17AP9PiAJh5D52+aznaRHsEdv+mf2vZ9+ZogkW
TQebYhZyWVqZeTWv+ix49g1joNv9Wu5OsNNB48Haas6mTEpHw2Sl1dpb2trjGOdp
FFHPCk5ZcQqn16XUKz8zAehkN6PlyWN3EcgvnpM0MHSYglqe/grjnpDyQyaceCAh
xFDmvoFKw2uPVGexTgFKPa074WvLE6TehGydRNPo43RymG+gtKsQ03Z6X8TsOVAE
KvAjNsiTTV81D5UxGaVIMDNuKEryt3LVKManUIaljto2QwFkZzgEljDbOc5BQJcZ
iHvc1/KDr7604dSSZt8KH+UJXn6hFN5TzrOPe9wS009SmMYHHCrjpffPDu/s11GL
KCkxlQRBk/YL6NEwqg7jJrHHEJsk3EdIfqKu0TpnUp4jGXP0YmUe148mOWf+XQQS
aMJWA/Q8TH4Y3tcUSBAH13xPgvc/Z8AEO9SPFELfCwX1nf2E0NWnjNrFtpzf/fU6
M04OPFT/JOSDqxym+OfE/fvxoCibMDnKRPFrlGdUvwIBAha5UHExrPk3kXeaYZ1f
g9HSxrwnZ7URzaUKIoJB0jszKmGveEnkPrbw/pW7E8BpVNkV4CxyX9by8YngHvh/
MGgcY5aiYV/u0vnV5DQ+E2LAt6P26829lC62ZD810jD5ZAr1kZTRXJJ6c3kW+4vE
uddU9yzyTwD8IaLkfUFJL9M4Dlu66iTIIzqwiNjGv3OqnP0YuLpWvn7GB3aifZ/d
n5pI35fgKOHrrqcpu/3/BwOV8gkVGvuotr4PDwFxnwzbqit9/glCk7ccy8mtucLj
+ovebUxav93w7ieOPwc6+k9kXfQw4iJV3rMVrwzkGiZVyOy6xWXctxplMcNlOEEP
F/cgs6sQ1fXv9a9kxiACFBhDNx2DVLQiBvg9fN4JKo3/0FjFvPTSHHsLx1R8/Naa
oap3lXztqtlJ/S58TNpv2QeKVGBP8GNLM9R4jB7JBXRoTSeiP9HsC3XwedCw5I75
hLUJzLpwkkcRFpvbQI8OLKY0gXOfanFEQkNboXQ0vdSxyDD+2mOIPUfKbrefpy71
uMavJH8voUVMFak146kqMGmTs4wmsT/E2S6O6qvQFbE6yzSo8GYJu9EukaVBrFBl
gvis7tcTT11HURgkKt7++hns1v5G9SVYfszGnVw2vTu4rvRWvhp/frazct5TBTrc
Ifp4VTAWGjZmtI78ThnRAMV6AuXCITv6QzP5U/joxT8B3NUXp+pb0CMLvOr1POXs
wwLwV7LBWE8mwxqcBJW58INJjsbk4wrvtrKFVStZ646rQdizqBlij7cjAC1JCWr4
NQpPzuI4pmFXXNYXBc4ZeyPhewUPax1ajm/tQonyaWn2cS5MKYEHvn/Wz4LV27NL
nPha9gTuyATc9EGr75NxGkHCUZ7MuOLwLyiKJdMatY1adUTAeTPxuA0iipfwx2Ec
xYQ2bpnc0jY3c/nNF3259i1Wkx6s1DyVoz6R4VaTFj8394asTfpJnjednIb1vVj6
2Avrjo33wwb+IXY5W9BNn5dB2ghxmXWhsO5OsGlS8qZXmb5Ykkn7QeWpzzyD6XMq
JXKoaoJYmoKWzkYAJUBbXV0Opeu1I0VlqgAXmi3O9Qs5FHqzyTgBm9clrpgCy1/4
lBVDcxuVrJzdXGGm6PiUHzHhxdGSiVZztWklV7PWtuM20LX8WpuFulDqsA0JoP/f
QEJHej5a+tck3sISvnf7IxZfmYSYaVp5RZ7VawmqXivywp+jQm2G9pzmQg3uCTUk
ppdOXx4Lw8RBz8SE3cUNfLH5/iGGkzjQTokCECzUYVMl/rGYUxqHFjwJ3Tn9kSF1
fz6LvOSBfIcPmSVUJiJCyp/3xs5UQCBoXYG2xnaXclHMX7vu5AYQiCQK2nNeQRsQ
KCTqbj5wLikP7j+tW5wKF5q73KrfafLVBcbYb1SBvN4gyxD2u+a7gIvm8VQFcQm3
E81bSh1fcLNRVBQLZphZhepnVqZZCUTnw5g6F7gCaauk2KNssII2Mozdzt0YPNYq
02k7rcwFK5Tj4QLV460vbUn1HZZQ8vCKyMiZvKRA1S6j6IUDFNnIWmg5uMgdlgfO
SLQA0oR0Jgp2B8Y1UJWUom7eJEIE8ykKTyc/7jkGFjAwYwGgqIZLTd5Ya7DAQnvD
ar7nVHTL3V2o6t0SFc895k7NQSeMIKccJs3gToHhNB9RKJqbEZJun+AIXEJpFTU7
PLu+3zcmMRlMm7wOS7t1n1HgnDigOrNsnmMq7hkaUFQAX+1HPcQVMjKJMbSTTvCN
3RPwpm7wPhpG6GoOjY/gguOvfuoP2aUGQfZzA8ZV2yLvj16kUkECJcvWZKUlANpC
peh4zHcl8olgA4S3S52aj0UzDyftuXLZzobmpiTNnoHxcz8eB2AirHUB6wpXBqKU
7DQxf6uNlLYaAIEdSZaa4sRAjUmu2La6SkNAK28Yhier1BMx95ZT49HdjzMAY2NK
pi0dl1Lo8l1OFCSs4l7oJKqqj0LTxHkSlTowBm5a32ruzcZ1kRiFvJFh0ZTkMNev
VbhG+wbp4BkDtgfoXVuKrkgR/yXrAtV3/V2W5O368Qfsu/RigjZFnWhQ8UmmpS2h
LrdqOVQdBdSSgQXfe745Y5eIeLhCKc07sPnv82iZ9/epe0bDkIIJPl42CWLqm9uE
wnHEVVAFFW5IS+UjTOCnGDmf93GpxXJEeOKzZvtutqI7B++2O/bhq0VNYAleMujz
RFg4EOli8lTEUNU1v9HYUSsiks0DIqZyul2lni/SZtZ8QQAf5qBvACQD5i6tHuK2
msqjaaIA0eR+MCF8gkUm/Izl9SDIBeR376OF3+Hn9z2lE7txzH5GM7j4tXHiVJSm
ZQPCreu+Ano+iNtYzv3y8ZE7QbXJxbPpa2rKCvXRTPEEs9a+qU78mVrbkcNdyqD3
m7AsiFnaFhsGqdrTg6K1BqpQPtpojlvMfhYHBgEfRPJ8cV6eU9A1K+bw4uOtb4NH
GXhs4Q3vbsrdHmidJXH3DN9ciAHEy6uHJ7DAKJUBtzh6JKk2byKXE0mFHWW4wS25
nKDNew3g3lvN2xITrnLE8OMPN9mjwiJRnkG3M4dQpdVrpkL5YGMrgVJlMI7zZnrm
IKsd+BB0luBKRxBkfnQpC+SRZ9vJqSO0cjw1jtpuimQDr9tDAjyUfBaNceYVPsGv
i8r/gQl5GEn4CNHeXgzt8KaKkaiQqxgrDCtEwzx7+6YdZCCKl2Bb/Fu/CHbOYvuq
n6txEzEyBIFd+9gPV+K0Pbok1KotDtUT/Gk7HuyUHRqQhaP1g8JfAcmfciVKp6nT
0Dt/EWx9zNPYynjlTANh9CkPJyK22SGg4DnVQh9lMyD/DPLmRobXB1dRs6CmHwMn
CDldkj3rEzpZ+KmwZFvqlF/h481o6Qd/Kk4/RIygt6vZJoinmNXVaqd6qa3ffpnN
o5F0WxvfZ+OSNnJcC+wxskMkgPgjHTqjpAe2I9gVurBbhBDQR3ovQreA9lHbPA8J
OErVjlCO48WoS+k6GSv9usO/NPGpl/nucR2xLbBDZlSW0vEVG9ec/z5nLdlVU1xj
Sx8qYH30wN2OdS++bidFDj76eH8cYgDF4fsFn4Z+jc79357tk5gwjsuU8Pztq4Hs
sOPxzEMcxHCBWTFtc7lcfjCgidb0Pzzg+wy1lC/uz9ETv3unsiOrU6K1a5+/mtOk
pyQWH/QRmcVIZnJIGClUtqKMywXEBkkqurxR9YcAA/z+oNa/17+diOVM/BKskDxY
Pz8rK/epfTHa0gOl2D8qj+IZMmlOXgyFSAGo0QsiNCrtq8vEwcqzV2si85h6Vr/9
8A7msvehi9Hc9G5TsX2JXMF0CFa+hk7amSHSSZzrk96JQrANnUW35FmykP+7yCvc
+UZTyKbgNLQ1zhktlhK4fY/J1liCqUxevcUzzW6cdW9mtjgtEaFPTY4mzcNvi3im
+AsAa1eIGklpJklhjbdb8AqffBLGvZvNOOoacKqSibY11ubL00fDYBkFdsCogeJy
PFgF3Wj/WLZx4g1MQ8LJRgBaejHdnMtSvZ6N3taxqIEJNjjrCIt1bLbPDDHX7DpU
7aScXIhQq41R8IyzoqFYXolqQiRYQzoQnoUYwpeuNucQjkXTYeHOYKiKQ1p57bHf
Apbaa0PktRa1xc7uNKYx5gYKlSBiet7Tp6zTW6BbPv0qISV6PSvIa81GC237BOVr
yXLjn21+KwG6ptD6V70Gx7O695tdxxhDwUwdyNkSQmvTuavtvbei5G633+aI8xHU
Df0QTcLNOwsL9xiw7p2VuLW7fP/QKhU32MdnMOFDhhbl9rD2OiPwhpUhIoGyHLGd
RElTazvSZf4SNp1EMsxtpGpYa7Rl5yxCyYJauECD6i4N1jcbLNAyKnLSjoMwrVbc
VOPG+75M97nDWW8naFmd/fJZpmumL7TuoCUSceTWx6L/PsEyXDrKrtNfqAodvJF0
9yfRZ6Iq5eoMwypyFveqZnSglPhrVUXzAnI2u/OWMYM9jyeE/TS4IGYORyXvdoHs
+pQ9om2Xf4EYFQM5v5HoTGyhS1ZUqQR0qNS1a9iLqneIsPPQzKU6nPD+88HPMgXX
0vWrGiZT9QwE/m5G4S36ErM4Ko41ObiYLpSDRZXR7H2UueVXZ3T6YmbhLmFM2Lnc
jdbJ7COrAp3P1uiD8l+HQW2zoKBr5KWj4B9ajmJzKahkxi/2Y4u4eWPDB9cI5zTk
57odqD6XNsmmUuPN9fb9t6UQs/8KarQNLY3aQ8LwnE69kKe3u06TtOnNHLNERyK3
BdVH00c/7XZEp4UCisS7oIPLOMK6G1R2aTRs4D6jfBSQvcRZfYpFerScqT8z+2cp
w7AH/17kzSVvZsL9IJ0jJoMg/gFiRq1kDx0fCcjm19Ua0r4M7+wRzNHKOYpY1ems
fud/ADqmdtnknqHbFQIsntAcnXJIO1wwnk40qrW2L1g2s8NDsE6brGD5AXZLUnA8
KglSZzPWTjIx9bjUm7W6MDG78x1sKTBLKjnNeb+qBzFQU40+jd++mpoJQ6UmLbLu
vl/0l7JrbeuQJ/kzIP5KeoG7/RESWVifmWPcDIjNkvNpARnuii7Rq4QiifkmpUG3
Hg9a+CWhA3WWeIeqjnCXuCQVy3FKsDqxlAVqz1RFGNPjjaYL5xYOUuwGB97hI4LP
q6Gw8BNhxOQ7aTSSfE6GWcofjovY/Ci+iHd6gBba1HsBCVLN3HmpPL1tYfIq8EvB
h82n17g1iFqOtxfJvNHuudThNn7k57UECt4jec4V0M4w5cdyPOzCuXLwl7K56lJh
ZqAR0sumD8w5NHiT5NwLibk3AQHJG5E6T2I5ZC7U3iR9WjnnjKgMDHAPBOa0i1i4
EQmqp8u1RaxTTNuSLkPl79DQPcegdzwDB+5Z2OBcNr7tm3dm9Vu+5kwQLnOXpdRL
KqvUAZQ7QEPEHF+pa+iG6aKUPaBesBlcW4+X7zObeK68b272w1vjd5zZPqDCwLhO
DmfRl0s+p0acZ9pNoDJMFIrMvzC9rY6zt0NyN805H1x9RoJiOd5KOnY2eZ+RuvSF
3Z6IFypzHpInHpBCnSL5VZs4FJBfaC7kJzIL8sON6vd9ne4tb0xrIagDO3lggnW3
VabvaRzGYq6+HvC+GLFp9RI24KI72OEtpld9c8DLK2ul2Eo8Hdx/jHXFiH10m1/L
lmwUKTXUpjlIXXxBHGOmwBMozp5+AwQn5PNQ/heL8+gAvHOcEda8akTOsn5NhmvO
VXww24tKxreVk3tMA2+r6lvpeMfapFwJsvFns+4VAYpv7G3FuKUoYxjpy7s3Sv2e
+7+4FBzG8tV9Yp5haBDC4Jg6mFeiAe11vr7PWTzJjiMM7BndiIveX+M6JWHhcArj
T9t4axNHZ65K9QPzEwcxjucP7SaN/HQmR50S+Z5S0vqngyrQqpl3CDTBzmKrpJWT
WaVOSLPBY745OfUcMA51y6Rn2lWbCD39wCuN46lP7h6L7Tj0Fbi/XPhYWN8K8chB
b4iv9xr5rtQaydbaqHsTyzEH8jDCvJDsteFADvyNlsUM1LtQbq+oWMFIu9rR0bBP
GlFSUA7XYjSEYUVVrE5gQ8GB3KeDS+LvSAUU9jSYcQY4Ct4HtKngOlUp2S2BkYkx
Da70hh7iEKDPWeZQK+OxqsrgoIg4dJLC3QP76aVnsyzzezRugwJuNkNvQpR7v6/r
vKQaSRoBuXToeI6CplaUcd5zneSeM6RYwWhPMTx/dIdUiUgtpVdVvc+4Y0TvFzIw
ltMhNKcwYA5j/LMX94pnHdPFKLxfB/bbbN1eVfq7neIpVJ2sOYVwpBupRB1mI8TL
4xfublJRxUsU61cYDpvwenM8bhYbJlqmNdhF69g03L5OfyTLnHEv8a8e4kK8Zy26
b8fTNh3ggxvsgTjNzhcIQQ3qdCyYqoIk1wmue4Z3TuUq+eJYFFyQGaJSsfyhaDK4
E8EmWw+NEmcATNv4RWEkda0mWRxxQVfz0DvFCZbrI+nh9nn1X/g6ndEyVRahk5CZ
8a7M52Rs2tFs+sAB0+LZAdfOIs7bqNCMclqaKu3pVIuNsHViONhpM6HGB+nFeogZ
g/DHY+yJKLzIsZM7rUmgKwCyn8c4TTQ5p67xE0FeUqnN+VIZq7s+AJYb0Khhp8cX
8c6YOh7N8Qfp8DIy4Dwej8/bjGLMl9+PEbPt4+4qctcwpAFVVzI+1tNJAcDTxscd
nnTI1FIkJlCi05JhstESGGsaPDtJeK6Q0nuQ/K5vJQ2BQeDNipRTypBOJT3EFMBc
Gpp+mFVBpLJ9a82eN15qA2xZ05b3XTgpbbH0w37OxwzSGlg5M4n3aGig9EYfBsOw
wtbGGUXnx7kqW3gkG74mPMxLmxHA3h6nSC2yVW+0SC9B0GkAmOGG9vu6Rho2R7QU
GNK6eXh17WNygd3EcxmaQs+PDUVIEKGl2uW5OiDkcoyCTBGZUu/H8ENUeu6fJFLD
iYM519vpQ+3mBZigJrAqfYKYguDz7GSvyR9TembZPY2yhSADpTW7IiPMiQN8u+ps
vfrvk1b7i8qgHJIdbeB3NLLtK3OiVpFiUjt7chHBnljvWvRUMWEVOEUEtLdvQEbb
6/vEpk5meNC7hfuHDCbYuDPicvqQqfTrmkZxhe5M3CDV5+XbhYCoBX2OATFbrks6
KdMlDRH+X8ZaBNwvd+dSRdfSSdeN9kyAE/yV3FtBS3WSZD8CmfJ4E91YF77Su30R
Yjn5aJZQyPhL5XbutvCSUdPjq7vMzQPEtrDCCX9ORSxFEFd2NUFt+3tJ9Dj1fSXr
HudQD67h2nlVtitfZTPt4e1m6IWj1DY7XAgt+ZJJaxI6dcDeSfG6EldW2eonNfmt
dKvhLZtEiNnxR47Y87qewKbg5i+jpjapIJIDrowBVptxW/Cn9ncXcLV35v8efsLN
ZzzMGDzFPerIO1vrdfwzi+9TUCSfh1Fm0J1LNmkxJfAD6v7L0F7djxSLqf2FVUC1
POSwmmWlkZ3qg0+Ti3y/IB3A963Rj8zEEcIJ+3LdmlsraSYRVUZmIECwQvemS4Qx
za35ulskNrcFcOq/S/rTA3j0J5N+eh99PcwkbZJMLF5ZlBkMYRhRZZez7F7h96Hs
inWiPTdtL2Gmud1LjmNJ2GRoJwobKpGo7pAmWQs5PB2qpD6j06aYYCdHqJopHWKj
1b1Gm/cc7hxnFVHNjUpoGA7ZvHRocgr7EaN8po8OsckDjmDFQizftT4EftLgDvZa
FlhhMgvtpM9N2aSDKryRfBL4VPFzvLA6YsA5OCE1KZ8mP51692DZrTa/IWKoGSaH
nwZRoD2JnsMiZJoPU+RpGOe3jH/y8zo59guCPF5KJKytj/L2/4CyhZkCK+UIgse7
TAm1SxWfc6RnuuB0p3z1qoMOQecAuaqk53isHxcUjg+/9TT8oJSIqBPadfm2nUTC
RBf4kfuwCJNLVkcYbnxaWBvaNeCEKPTwESYGl2jtwHmtV5Yt9C8gkj4MFPXubAgN
EomNqXVcUp/CLPfA7dLZ1RYNYQ+pxPSruAG/JShUWBQl/dJKg9D5EO9Uv4PXODzB
RlWQjGGEXFN6DoM0CPTJ1PXmCUIYOEdjarDmEdXQa+dHAJTpWk2bKY6XUgwOWRwC
i756pqczSSY/5jEx56JzB8tkMCGc3SP+YGLmmr+NXveeSHfLKsm6CdXfy8/tk+X2
cFpyasAjJtWBNyM5+166jgDIzZrfM/1lqpmhr/tTWvnTNsPFED6RMLwziFpbjFsP
z2kiBVaHeQ6+ju8bcYDXjqHwIMMXAP2AI5/bBnluJlBysC9As2IMe3rrvNfzEYTp
FC504VP238v7t4rhUTyIWJt71dk5BraL2HzX+yRj6GI741gph+JxKL3PBwTf9xeb
AbtRzzB1aO9iH00UgzRLseHYvoD5BLmS844QcAue8tfme0BzjmZeiWxXUwCUMNTt
Z+xGOF9YgIFIH2Kff/47OLXtgOWMMHiLlZheMpNpz9/jGfUJp0DtMRWL9jIFCajS
+aEjYbH+3PS339PrVqXWYKYdXQzuyhhJ4E+3GNhZCRZ7nLki6mi76rYIONfB2lJz
GrWcEq1Q9dKsj/mJRhoPWpFId79J44KASf6yDpb6/p6ojbsY5eItKQpsJ/efgOLy
Kt2Qi08N2ZtuliP6gdLn+zkExCOcRlMqe22jYsw1Ga6tq/Z6idpZ8wFfSyigeX54
jmvJhL86qXV+9dTkwLpeoak+fsXp5ZOTDncveQCR7nVDy3A5OOU6sNNcK9QKm/3Y
svZcUl2kxQUH4nAAnvRG6vuPRmXsHJi2wk6B7crlkTj0h6qdPVbcwA/ks04fGQXy
yv3A7tDcH1kR4F6pYZ0kQjjkr/ZQaXjwd/GWAu2l0IQnRvXbNSJgiHnpNlS7YohO
YhinBXfNsJhU684RehKoJBL4YM0jS2Q47sxgEeb0UUY1Iapb8hwYJAcpolWY5asQ
QsZbN06WtGh65h4PNPCiKNwm6XE1tm/q0Ubn3bxQJLuD0Dyo7jnCpldEe1nm5tAl
UBzr6VcHcx+zcqz7FHT955dJE9rN1cwRZQBPgNMWTZl/v99uso96BsEI6JpywB1l
y7moblMkhCfFCtmGK1WofgZVIirxzqQvfb3wWXvlUwbCA6o1l8F9FMoBc57egnZG
IYX2nR2qtuTOGlOOHjRpwDphQfs2ntDLZS6YNs+eeh+Y3LMvE4mGszT6Ms/F2MjO
Fsv+GzHGPtYLlDTMznrjtqdMtj3sAYBs3hgaX7bTr0ml4bjaFWAkFmez7Z6Psgxd
eqJKVtFwoC0ANKmIeNnmzQ5HMAZjl8A7Qb/sCObi61kZUF6s8vBmfRXGWnewdaSv
B3HsKp/v8vvGTVzf6T2ZYhO8ijGxWu2RUUFLldduotKjJ23lp5x1PLh+SccTxI32
BTlqPv2d3ix69goHbOARfFFZmB5XFEgphB3/mGfoxI17zcrB5Xisppp+1daMk5kk
r1uaY6qo8X8MpAbXSD0GkIuZwKhRfnbcwa2nQLJ5KKVTQgfIQZLSFQkY491rVJL5
pCiS+NQiK7/y3Tu4rGsk65HHGXg1GGXYjjnk1ijSaAYRCYmgkZ00petYB8qQ8WN1
iGn7EL6J+LnQFsEfl/hvtBgVtlVyiEUIY6cTX+JoB2RdvZUDk8tuoJXA3BxjYnEU
2EKRKp8SBEhPqA1DbfB/dTYLr0rQSFeGEgWkAuGz3fXTke/7OR5tXeTuSZvs8vgk
XAurs1Mh89RB63/SgKqu8q4EZ8mFDr1utgQgknKOJO8+psTT0sCMXDDV97qwlE2N
ZuoZGdosiLv02oygL4xlGI62ucNHsMorcIHUxNVfVWbY4+j79CgotaJiEsfKKEb4
qRVlLi+T3raij3iMa7iqjRjQ3I3m0GYs87l1VeB5iwYWgnswUCYwDR9OZo8MgRDc
gOLzP0KBi14nD+39yWq4CwsnSzz8DXA4VKCe+6gyqVv9Nrmik5wCxzGG3BAjTPWW
2l6IC4LR/gK4HWJTYwXswUQJBRzuUm4PpX9L3CcJ4XncStasKzGmT6Hq/MYZYU8n
zdzkaKNfA6nPq/tgBT0ySBkRuJRxXsIxFOeaIhVn+/E+70sRBStOAxwlo7dQGGz0
waT+dPkAldrgC7Cha5TXsFsbiGxCvLzfWSrDoniomqZFb5WSltESd9mofIqw4fZA
fYTZYbX6XFx8suHx9eYZBT4OB8XgniumhggbBVOkM8actpotoZ+yFuaR7RH/CWBY
rKp4ca8Sxe+yMpqvUYFG/RRyGlV7K5WGKGeKCbQIP7wgH8GQj3wBPiGMsLHYbw+q
GBXC5AiHS6BhKYhYzCI8542PlIRCaYIQT29wOh/CjbJdqXMlJ88NizW6zAl3J+EI
JQVGcTN0ScEEPwFcvOF+6IrfG0R64FXg+DhUsyHl1K7UFI42OJzwf4gbTLs1LJR7
UKZAEQIGA3MsrWNXisSiUFW2P5nuRUFEnymjtpz02K0hbj4SdsHGv9Fl1hX2+yQU
Rmon0ipW/wqPCRj7IrNprk+oZuRaEItsoS+zpbgUR39fE3UzmzgpmSD35slKsu8+
MlsfkCpz3bUlkGVXDGsY7OSfEMrq+s1N0l2wi5S2UlkCjRs6RqnXqI4gDn7IvF7w
Rl5pr7KNoUewj1FkS8+QT1iswDTS9F4nCQu19LmEXKXJXf5RcZFUL+eaUosj51hM
IKVtatWFOtn+x80VzJpgy+aYB45GyPScnPMMsVupivcbRSZayONe8arH+rymWN2s
C0Yvf/voJMYF85hmhW4BG656QKlssxgzhgy588ZWKHbedAmTJEBOhzxgsoUOshbe
93ATofoSdDXESPezRWG0H81H66LoxFX7bD4neXPdpZN7aWUzzOAhhpZrF8e43lya
06bgXw/P05D59ijEQw5y493wSQX1EnBJA8Dba/J58RF4LPMdyvag3zQYXeLXHNeJ
vw7Ef0AnCxG0w11EMfYmyra+aPWGPTZ3KVvfim4QwFuMVdixg8ZQ0OLwXm5MQ/0A
cvgIAo8zAUBs/LM2bVW0Is0VaqS6Me/VOvYygW1IxkfVgJ47nhgvcH2rEvDcjGew
iQyxFIQmQl1qo2aE4k3dn6HLcbmoTjD6G87Gbu9WRhIaL7p+9odd66CrG1jlSjhA
Uqco1OvrcDEMt69otfk8wpOZBcTfmMWQsnu/nwHeUYaspLBIGPLOkTGBStSSuIdu
OiviAR9yGzK0SNe8E0JTi6BN17lXSUhc2zmzEn/a1g2TGq7tiDm4hRvArboRmmnI
jW78aTPNxwdKM23FZLYa8QkZr49KiuUruc1i1rLZHOsqREUJMMz92ELoNQX0od0e
gHCmJkklzhPGMss8Gz1UkaQ6Bx7mVyApZrtVJYeK8pfH5ZuPQpO3BJiYWAv+GJor
1ner2ZfpNo1HOxf5V8UH5vassgR9BlGZlJAlaERR8q245wZjKHlcnj1FZqbPMZ8W
X68FDNldcd/MbolOU4afFjoSHsY70enVGth/cTb77mUixAOfrE5mKa2/U6uiyCKw
wg2MCiXKefc0Y5Vk8nBeMLXqz8F52O+DFy1BYxMm+0AYE9pydVfwtltENOBoQ43G
o+HlZWThkAo2joiMW+QMEAiGFnIcJev5yu2LkJRLJl/Q1lNNYplvE26J/S5ppBSn
58Ea+O9jv96pP54sPi1gdPb6skyuPLADqm0lZcIUScW5ThfIYWKRuMT7JQtoH2/d
a3P919AwSn9DYUQEDeGYDNNbwwiHM29BDUktAzSBbg4ZarvpLqLIpc09FSR2kdGG
pRY3F3yP66DIvn43vWtGpxCkp3eKJkviljwConIl7eeh9HZ07tyEoO2AK0oVok2E
NDNzQFqiA/RvxZyLJD2P14d5OU4zylG+FpuokV9yc39sPVD9s53ZYSWCVmMqmZqz
LLq/GFC5xm7VdTkZHDjJh2/Ah66KCoacJqZGpsgeP5U028kObwlvSC+iGaEHB4OM
kX2/PXj04H2Cip4un83dDhzX6V3nKB0iQHozRIbSm/8cs1lNAvrpXjSo9dHN6cR9
1OtlBxoU441InXa1QDLODCgM6E/dGK5W2q813Kh//y1AmIC23iPWk2RLlGYNR+4u
rvu18sd8x7XTxnGrKBucv6GfO3jLiJoUUgA+TeOP3UlvrF/85WvjhZyClL9cUf7t
7JtfmesWMiXfcL3Ax75pPWVN9UzEbDhMj8BXGqTxo0CBzZa52pLTRAT7tDPPvVOc
J7AOPDV/3X7Hjt8QOQGNPk1m9O8YmkZjJh7HGLkhx0FXNn7VWY2JWi9hewRy1LFc
MKU162v08GGOKq9UrweKE1aKxG0yw2oHwf48LBNyBa7ZMWUH09lHCa779RcvTghb
W5DB93rrS6GkOC3/fhN0gpgkaR0F/DjO7/kdSs15ULqLxUE/7KiuOsvus493Cmx6
oJVUekDbK8sKKM+ijqlQGwiOPgLi40hbsse3D9tZWbG60Q1dB/cM+ghJcydvHv14
DI4XWgLYHK/mB/1wVimuPFk+XNfe2U7ktMvGVjdJ4eNy2zUCqu2eG9usB2++BsBu
ZOdxCvyc+jcFZ5qDs4rCeYRBUM7XFbdxEwC1S4HuE1VS6beC9VZEkjmFclPJNjws
1vmo9sTY3pdCt8JrQ7SuBJ0bKEGL+LVP95uMvQxXd6jwRueLOZ5oPO4p+c/k5yO3
3XGXdHo+stoOV3v7KCNwqxUNeUpu2jBaNeKl+uW8ddedAf79aIz6KbfR6KYhkfMl
bXuZzzC2xWhy7zDyw4IfgsYmRb74Z38qZwQZjY1hE0aBvUyPdvKDUPZjgjFbFUzY
uRDIpGWEc+aHcgCsVOWtTXytHE1DGokHtPYDDmcf5so2RY40WFxuA/EVu2Ub7aCb
O9M87YQ+GMF0FEp1BFOyZ7CKacknrqL4tX6eicdM/AUMbADLvMygp72bcOj3nUPg
1zlSOmnasVa3a1lkHbabk5r6qE3bchzosZ2sSkuBn3CxCybOqTuZjKJAD8Ja54A8
+JdfEtKPmRgUtaBOxLymxb5RHyNkALqx+QRiEY9RkboiYRmF8XRc10QaY0KKpBt4
3Dv5GPzxy7v783++MXtfdd5uEvn5s3NaVzxX64QeexgXK22SNp+PP3r/x1sCASuL
HL++AGTfe5UvBS9qHabMfxeO5Cf6pv6dQzyUH4S+9NqVy6SbOTVFZkZrkaahLrL7
WHd1sC5o29CMWCpzQ4tG/5TsPPci32s/dq46BOTCIQRMBMobENeDK4TLe1TKvUyn
NIAhXJ5rO9YTdeUQWg/rNPfLG0V2IfUadrEggT90oJl88hBzPdY/yeKp2+acwoTZ
+W2X7b8dwtLbDwe3+nFTnQykRQH/aUQWfcSV4ti6RgAaOGGSkhbmmK2h8NQv4O39
lN/Mhl3Ltm7Y5D+XvIJWdxJhDMA7tuM5A6WWODIF3+fh6VvB+1PD2HGDaCDGB9U1
boy0myhM+ENoqmlCsVILXxWhPe0lxvKjutigvMecFO1hooVP5c5w+kc4vhR/NO3Y
y0ItkmQa6M/ppIjsSRvTH6WHlfLEVpNiK41wPj8Gr6O1P+05YOcnEDs0WJq1D2ad
U+DI2gdF0sf+YTQryyscNxdL/SDqBXF2FCCtuLyfFnKdGhl2bVxV4A74ukCkHU91
sfVXKJH93Xh/z2whbmTczTg58s21lVsjd+D6zTuPBJL4naz+7cYCm/THGE8ulNWu
XPHb60gXKfBsezXSpkCDvso+fyvmsBmlBz+GhcczhpPooNOW0PSyvCaUywRKqnFX
9Em1GLM2j+agrqShOqpHJ8XrmZDefJoVDNsvujiQSjDcd8Yb301H45njhW4NFI0i
9Zujjji78srwYM8LYLBUO954eIykoOEtNw8qfZ5P01Gu/MM89NkT6bBrGxuY8dxn
gQf14wUAaDTMw2EAf27pzBnw79WnYWkzxXoxkE17rp7vr4twbENrESk6/dYTnH06
DU4sAGPfrnh2bwN0xXbi4IaOLT1sRy0JPP/THok8qNiej3uTDDMeoJuEdPAy6bUg
lVAyQFNRCAq3Qj8zY7BjsbRPRjNFousFnw6R0IO6OcCRkRg9eV97JSOaBGloOAiy
agBnkBWq0DTigI/uJdUnygzSwufblvi8ysDYXdZQw11tByiM52E028+7rDCQH5ma
KefF0Yf/dGLdFRk4E0v3YRdebN+x7Z6uE1AMlUeTuAuyJJYQRgP8jchpKp3DR8Nf
0TyHm1JmxNir8J86jLLTJFpd9Tq6LOwm6NlqN2FEuJtpoM5EmuIyViFD3SGi51Kd
7Em0gs52vxHDaEhpTGc3xb4DiPlVb26OJ4VKQlHba1pO1QNMhoK4noGHPsAnUtWx
yFEVnpWwKtFaVzMHPIy6qtudNYk4b223T9Z4V28fcVUvZxjQMEGgBS6CDr7i5wBp
xDkWAOffhtm8157zfexyvwl+DhBwCkZhM3HBbhuu8vtyYHHmraxQ3vGGPLNpjfER
bQH8umiPC+jcqoNbEEskdHslT0LyUwQd2pyXRUtzMIcZMqo1w2ZIw5dqIs66Hyq8
el69kahLswFo6KW4dqDp5WGfi42GGJwtIgCHfyNd9IRvy2FUJIjbdFDjOjp7ybrL
TChgLtCBXbIBljDnKCRQcihznqSHvg+4Y5nZfNVYmrhzHpQZUJwt18Swnh2gnwIY
gdwaKuflmzI2olPWZ1zOqVWoVrn0I7gY2DshZ2UK2tDvQcG/O/h0dUpeXEpQsGeS
+9nlhFzJ+jGrukBs8DUEanZa1Qb6f/eAVVU5TDpYSt158bsvP/+skSwWeN2IkDXy
MGGxb3iVLXzuMybM7JP6VyLXQhtj1Wr4I18H7m6rB+CSSLH6s3FOaLgO5tiSKJfp
bUoZInu4TaijLg9gZRrATsrN66nWKRkNY3AO/+mMXApO1J0b3NBIYtFOfnvXjX5u
MrRZEjh45lnNOsvtPajp1XCd31C6mSrCjgSA4U8pzO75cSvhmEDn+NTZo+Njs1QP
VQphAvVw1QZ6PZk2vZ+4W0OqrDRA1dauqIOJk0Bi9nubskMf3oR6Q1ShmHM9wr6h
ksy20YrO0SEKL+IM0fWloLzgDSLY1p6XSMVW4DtCkPVnAr+yri7sZd/m3qi9RcTF
cPsdNJdVsIYXyPidMGK8A94sroWfKJrg+GrIMwVSZ+kcZwxPy9RnD6B6lw+VzrTJ
WTh4+o4oJeCOny94tZYwrWJjQAkWZMHXG1JvLkoiVomx9FYeKGAoV3cBz3ArYq75
QpuDXOjcdD2GQhBohtaIAs18uK7gQEqCRazXYyM947stwBMGk2d8AtbW6Ub0CTpm
wzmwWZJNQg0ZU8t1Dp/OjJNI5QBohOFoN3RHJYEB9rD/MGsML8zx3oOEXEcUhXOS
BRVsckuXXZTiY85dWTcY9raUXLLZKy/Qytl6BGY+LbVhV11K5Vqs/wVMK4rSkRpy
N3bEv6idzy6PtRVi+03E8nWugTUSou9gChGET6+MNG7XQLMd+lPX9OqZiSIeoiMD
KiKUiFMYzUXCTJwWPGQ85vkXWv8WvZlFHN+VVoy5xpR5Cmu5P4m6HOcPIeZf0KEr
p4gPEQGynNzUQyNFrCxzrmC+Esn69o0Swt9UhQ6eGJ9bSz8rznJelbZF7qWNN/Nd
utWEu8X4t1JWLPzCtfDZ8pJFcGi2IACTFELrG+5x0NIOeEzpyLTXwNRFY/JmnmAs
QtLpBkfwujZMpyePS7KwnZmGOvIHCFgZQO3Yu8oii9OviAWJz17cux9/+izzecmQ
gJOPZGco6Oe/iojNlteHEiDKJloWAwukatHiM1Sw0mDBLH4M0CuSje/ZKhxjSvRY
SYQvLvpEhTdQDaCubkizrnKmnTVkpBg1vSrzG6qsGgz3NQBSh/Dzk4dIqlbc6cb5
DTE7w1FjSLHy6Gg341S/2agrSCRLKcQ5z6R6NVv2HMv7v0uCGfFKGVLaXZpNtz33
AsrsLp/5fV879MnoxMhZZPt2YcxdxpN5d/FIJw/ukATlZkVzeXgD2RMroHBuvCe7
L67fGJM6l7RLwekYXvh48thIYXW1bt9fKwztGhW4P0vJy8GgbyyldTjDgpwmIDMe
f72u+joZtCztMY2OOG95eV3yRj6Kd7+Q9kAQbTA8iWiEzCtI94YvqlzVRiIDM26C
K7kD/iRX4zAyBKnyJdSxYyvIN1PABmu/boy/Q9LwVP5JCFEWmDEVNqY8hjtS6cv6
y5iGaW7aBv3HOa3/wvXrfdjEU4jB2Z/JPXuRLAWy+cJBn+NU5txTV9RQ+u3rtWP1
ejEFiDnhUVWeza+svqUSZcTXybKOCc55NDhaLRIoaK1ukJJXL/z8Sc5reHFBhLta
TxeFhRAPtTnSrQLdJupUkMLOhrAe8vCz8+6o1Q2S7StxzcFaVtKQFifkKZ3RdzZ8
FZZQReXrgMVgD0vOD447fD8lA73/ffHBkiCyzj3PhThL2fjYPhc/3dsa9OnDrhHt
ur0PCe6OOiyoYIOToJpWyoFOgw3HmcGKfgEAjx9syXKsr6zNcPn+1xnn9s16kvtr
r+epqSKciTMO+xuIaxvsBXlTzPZqY7raUO7awF7RZSxUvcXM7VZCyoorJtchcymE
NC4S5geFocq/qT2qtaEtUGrx4qF9rDtj15XtfuwFl4FtqT/mzBvyRsbYeBG8gqpl
qUcyuZZBdkt7GiRKvW+ohAwrNMIBE3IMEs1Gx4rtfAAPifQIsQj/0qdis+7pblox
oXTld0g8XBLkXo+YCeGo0OFg7towNFc8I1yAF3ZiqeMxGoteMd1yJdl46DtcYPRh
S7ByUjN6ELImZAK4mVvmSznr5cZCkLuNhFjXZ2s7A6t6AdeWinqHPxqShGGuZ6nY
CNaxZnCrafOIDRB0b50W5gNNf6q+WWQ/00+5Z9juGrZdU27qtEd8wD8FJ2hSgExX
ZLFumjcS/uDhfmgj55Aj6KgIqqqaWucK3+qnpB494g/DMKHq1TugM8aStSXReKBI
E6auHMpZSvmiJ6mU+UxxYrDmE0AxfhI0gitTY3BOhTox8Baayj9QnzO8etSSsZZg
Tq3Dkux0rgk7juWyNNKIeHwm9KSGRlEDbAXhxYDomDT5fw/GQwidqj5FV3/71ZS5
vACrcc51K+NBViPQRutkQgBrMvagw5TDLWNe1DwJvaYkPrKa8VPqjyzvmB1pI8F1
JuXwYjoI4ageU0N1WqEM6xw9wRFGCzzvtdRcHaPYGbbobOjFA7OmBRxAzapIw69Y
R87JfcU21JowaGLz4KlplMkg3JpZvN8KMvexjXdP79MSczcOsT4ZIeWibg3Dc1V/
tspjph+Sr9Sv/umlixnQWR2+tezSAKDj9ZGXQ5BCX9zDM76CrbxOGR08JuuCPF+Z
cPdOOFO9tR4nSr1l43IxmZ3HMu7nL6QcQhAWIW/W8ySl6ZdWH3qZiY3dpadVBMme
814WLEJqlvVlPWZZwiBonY4QeObu+LVKqkPYBdTBh4SywmF6bjUjlCvnm8Ub28kM
+sFvMLKapPykoiLjCTL4tPsp28BWgglGx1W57uvNJifwolQ0qY/LxasSfcWyueDZ
AYiyaGpqRAvFdMkqZ29LM/kvtBdCwDrRypwky5lQv25zXHcA5SVLt5/2ijrQfpH+
lqe8Qb0D6G49wRzvySUffwcBy1gcfquRF0hgelUku0n5lxTqujZOg0Np+qlbm3F1
ta99Hor6/kapD23e4TQDwQfAI0GtkYQ/H5HwiEnLSOpS00WQUM1TevIKpz5To7iJ
NXQshNi6Ow0/2zQXgdNTGOzaca+FoNUD0AoaR63UrXv6yNGPBlcsrN0/90NESmIQ
tctNlVJVRzw16MjGXWZbj7EAJAQ1DmYNqcBXQSkld6TGcKlx+GDkiChZNt9GrulA
13TbeEVpkZAnCG5LoKO7wpKGoH7cQxI7lHCP/Am46EXxx/OrPptkcEMLCz7kLJ5o
sOYYAcJdM2uus2LCg28r+OHLHQr1BdbIXeEdUqebLASU3WJyjeua+35FS6zrsdTz
JOipTahXo9ucqhNyCo2tAR3whc8Mn4WJs4gwYbSgcOvvlZwW+sY9oLwfI9j7ikez
s+FwYm5OyEeKjuFiGopUc1C1ksFmGMzNfGsGr9NVPK3O6DnK2HD0QA/swCMY6AIu
31RLc/ro1nPKse4D5BG09q00JmyZ6dZUxpSOGQG4emsqx8+LqHe6ocZ+PZgs930k
mQr+Wof6P6g1KRG/GcL/wliBgzD7BLDIuHMI1MRezo9H0Djal25UzpaPsalNz9OJ
6azTjwK8u5UigxoDvq5afE0w0QAqTEyYuKAQS2OyZGElPvdHK7zgiM7cdPyr64dW
Z3PZLJWm6N0ChWb1sFQ7jXeveJrh8Jpy+Y0R5yv4Z79LiuVTz8mW1OJQkcS4XPOZ
ikqTz09k8feF8dyB4DXM8RaUEWl4Otwis03Vg6izSHckW0fwr1ZArh9gDQWbZg1M
94zryG/jUBc/PK0eX2yuspDVOU9p8C2PPXpt20lsafHGf6nrDiqhTELyg3yZKJI4
zRgSrJ+F3VT7Ee71YrSl/ISKhw+d/Jwh4/ENtghLnF1+D9cAVQRQk2YPSTdy0pYc
0GvbhKuVrrvzLaXa9iTDZx77SdePsB443fkKCP8lSDEcNbFBOk7Lh2xkEdWf5rzD
mpvc6Ro9vk0SfR1omUJzc/XeiNClu6o5GWw96SiRy3oeCtCNCmF7K10bLp1XJ6mU
jyqFP/lgWgQK7mzrHYqrZoVmQM8ZLzBMWQnXT1QrMK7yFbnh18I+wo82WcA8+WCl
dDw9b7+an3yI6ixr59YDV6YWs2MdIneuObYeHEqk/Pei6/hS5KXy2uQoGaapcpw0
hAc1B2IgE5tx1hHtJOHBrfhA03+StZRkjXZn3o/8GFLYJ+eTJjRoypoZUamWbj7Y
TTqshnKtm5koc9dNrURfbbHJIISAU0NTCr9kAMfkLG3mw9DdLm9eZrXQMav+Tblf
g6nwvuolMfM3apG+95JmyedtVzjwTK8nf4AQC5YSMU+aTsmYgehj1DC3AI8mnWET
Hh6Bi8v9/nvdm1vvbFXb+uewmyNnWNMCch58JN5rOvgi+zyNq5xmCHfB/w8qpDJ+
ptZ+odjFNRM4ohNqduCM0Ald45wWGCODZm7dMJQGKU5PYst2YSwf8dqOoo6SwqPn
h8BuVVh6bf+4P49lA68kXGN5bjTZr3Y1nh+XJlvUsCS76Q8AEhTckczaGVceI4zx
BnhW5zjg8BnHB6N8WAxF00vnzMZ5qcomvvG4ELW8Ad8L9vYRRXcdwwfN/XGBQPAe
WqP0SV+U5UGlrFQi60WBkuYFv1iw8Bp46NRwIGiYSPBLYETV4F/CB/+k/+mZ3/ME
2gzKhZ/Ny6jHVuv+M7Rm9/SL/UTwvKuIsfbOL1J0D/1ktLhKzyFrEBA3ymHeMppz
xSbzPxy4VJ6ynrwHMnsWRV3+x6Fo9Kcm7sepni3T5dcd9VbN+OLLoaGh6RO4gLYM
1J1JsZG9Rqp22XOU/Kfz7IPV0hTGh5Rj+YlE4YCZxahUagfZkeOkfOtABjESU9H3
RfA/gX98+qewqZPkZfr5F1YDdx868SIsbVaUh/6i+jrcHIi8o2qjUksfACjRdsBP
ZUb07XV5jeh5p8XAfx2RGy12Of9dW9XDcAm+gqbVXiGIwf/9aNPy9IrR6dpks3cS
LzzDGGGYfL/aCjOB8B1GrPvb1iqUi993nxvGBxUT61ud92hNx7nosVPMGh/gds2M
cnRo5m4Qah7/g1JNNkm0hyNk7UBZ9XrhRI4A8wzb4oSAYKUeOH1+0g5Ca4uuAcfw
FMekoOPxuQ/86A+iLetE8lqdWeRG1Fss9yloSLKZo+RJA9mhJkrQKepgc98fkjsc
79c4MF8Kf3hyBnGR2fS/8MaE34dWAlZg7WLCK97iVu9Rw0kRJv3WCz3DAK4FzDx7
qHxZna5ctyEiNpsnmlc1suBj/bDyTGPX1x6yevRJzNdohsZcYcRI5NlG5VaDlz6E
EOxK8wLm1MN5bztSo2pzsz/uDm6T4iBajT1fHriAIAS+L1eYx0NBYc7uHUb+hEEu
DfObfwkByBO8czYN+h5kYO1wKiI4JUiKU1AaDPyX5c1r7TGRw4s7R/LFKSC3JTsO
3TZqBIXQ5+gnp1PkAxTF5j4OzuWxfX/u7quo0z1XWWKCwbPkX5ztTgkTzJyg24TN
N6RIqo+goZiqqOFaKTozqeIxNzN4Cu6gICN44hwO1hJ3Ca00O1Ln9jEhQA95PDjZ
2TlQzymTfF+xaceJ1U7GDIB/duJ84zOHMIyH1QEn9N+5FzrGfcdObX3rLw2dLusm
NpYDtlwLEua4xsafNNr5i7HnGO0BfOSGfqwWmO5nR42v9MzKN5VF3nwuXPu7JKVj
8hKImTg+qcZC7C5cjpsxxMNuDRUXWHDKYQRP14xpRzzQYCGIntT5lzx1hZ4B/CbB
YJk5wIga71U68t3BhjfODprBhAEGOUWiKST1J09V8WQZyLIvg6djKTNf0sMZk7Nr
JGg2o2gy1HifQ7Dnie3QNn2cj+zczYSiDysU2soIxSuC+j5E4PxoJkk+PIvR5sGX
ZJky5SBb3IHjVl43LJZR/HUtlfflBkiy9MENaxJ+dxmeS7Mpd67+xVbb72syq34w
larC3V+a7CiPqw+QgmgjP1cnwlLfQjFdylMDM/R5TbIw6hDdoKI9rW4i3xyXQN9q
8S2l7n0XpW0VceTZx8NqFyYZRweH0J8l7HELao2B10v+kdho5CgYa9I0dVDcaj20
U9qAjEKFmLdyHFHkeVCmbXJb9aVR9DXhut5PqrLRNTk7t/dWmKGvE0qaMXlyFKMb
qFq0NEdNXjA2VWGboW+pU9XBKb3ApVlq9soOeo9Zf/x9C+lrWYa9P6hPOv87ZfOS
Xmc6qFU9jsNNxHkv6cEGLEiac2WKiLf1U6/SPlJmPoQRcQgChgFWRF4Wpb4grtzU
yMxpMzB9N+I7l+pmwQ/FpKoXrWqiQZBrtOwy/KWDvjwf4X5eQek3FnUYnxCDIj4j
DDjHtYuXojcW6r3vjsmN6wjW3O9D/imeY/aAmvO/fHFAq5m8N68ae+rhBf6rSKGs
yAoSlrvUNrGVerUG8JcOo4gYwz1kW6Vy1yf/UgM9sKDl45EzsWNiFVk29WlLkb63
FlcZiNOBABfXHuOyEPmF15stkopXPJaQm9PseAD20RUMXCBwgaBYLVxaDtkgneyV
0BAoBz5nqxgggEO1m1HD7xnOBEs1qZukNW+fL0D1fa46nxHFzQmOqpzwvAQLS88q
/ZjM6tbfd6PHaQmuAKlWwj8Qo/6iLwn17nnYzStFHaasReL3USxNemwfxf3F9L1y
Nw29Gbv5qD7h8HKp1rO2ojgGFO37lFRh8F8rUAcm8tRXDk85t1BX1RKJfjtXcFfW
QzuBTTcT2Uc+8TEEZyrZmm2RBbzWAVGhGbLhFf5tpn05arSV2vJKR64hJ2Ta2QjA
IW82uCjdJovHIwEv0LdxxCK3E+EbijfsehPsed0CY0/OoBRzGBGJNHxYqtMk6I4U
lo/iADo+aJa29MGF2l1douVd4CZnS11MNYhidZwMQYzpFC/PDE9nO4Ts4p+PcRXH
eSpt3qa2Ct2PGUrObUPPx/GzcFFsDqEeKycPJ1mH5quEwcVvwMqTn/4PqPFOBI7A
VTVU37tmOMaE8KQ3E4hcyhrWkQp0MJcUCOyImf9UIZsFPSRJUTCKhZi2uhtA4sar
7+NgBsGPBFM1yZgFF9+ueVORPCFXi+Zb4B92/3BgS5z+H3bBTAEM9SQV85JlZICM
/osihGULTl6984m2gRSF4Ijg/nZ9m8290ps3ryae523YQzgTIseEtweMZZq7RkVD
aUc567gC2jSMctJBa/pi1xJsXrTjb5ZeY6WiZSN5wrSq+kbIX7/4viL9CPdIqEJC
51B4rzKcHE1y4qV8kY0uQO4Gsg+0FnPKDCexFIP1C6Zmm0c23TsTbWPTS/mgd7xm
C/mxfbOQ/BlHchrH5WGBmik9jWUwH+kzciVE+YhTD/yhQbna5R/LsSR7izoTNNm/
2Snl34f6HHHoSPzgic5+XDWGGEsnDX8WK+DpSkEDro/5kQUMdk5DiZTc+sh+jYR+
+ldzmEhTRKcxjmgygDHypfZMUm/3Cs91BIJTRMTuEckHcn7Egq4c+562G8Yz3XZl
g3Bpj9VI78fJfB5ns3h2mPrYGEQAYNwlSC55JpX5lsQqEoCfUT+/JpzvtirrnJiG
UaJePBz7w6XQ/19CTjKdEhdgmtKo/+UjTDrxVpOltfcV5USEO7ZOl71SMJN1Oqq6
4AjJLmXXFdDGRroV5jeop3pjjW3Tda9GRt0o/ebAOaV1yxglzSZmo0WZPhK1WcvG
s7n6pBHEC+OGbT3GZgPvI1TE+ezPeTS2piTvl0N/9ArkDyaDlS5E0yoq4wdx2uzm
qL06KR6TAKew2kOwU0fMfHe6fN4kil5Relm6FW2bvyuPI97V1NcEecGKPWgWEyMO
BkmLpH826aEnTqYZwT37GobhBJCpKu3rDDyvsyXg/O26ZUPdQXhLDDQ8FKKwmVAL
tK7udMrydCUpeHB/hKvCEowb+NyocRKRDsiZsAroOXSQcyht4MemrPxjwARTGBOQ
HF4U8haVbkAVWfLjM2z8m9dlSi5jQuvShhosJO4vGk4ncEMQKLPRDSKFY+oGCy+z
vt6kHe12RQrcqH6Q6KlsaePzBmt1aCat2iaW6BHJntBbCI5AvnIZeBXNKufWr9lz
1arxNoToRheiadSFVF3ywaNvnTaTFqnAwSD8adtnL8RhGb4OAFCT6JaTrVVv9f9x
`pragma protect end_protected
