// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:45 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WaJwXlLiw8VvgDvgvxA4wZbowKI4qXZHSBUb898WY30xOkX8ZUMDkUY19Zc3rAh4
ve5eUtZVSfbQqOLjdXetuqiEyiZZtLEROzWP9qsEhHn1jf7tzUxbySnOSaJejDYr
LHbmjPKT+4/7A3unfq7gM8MkEr9izt9J8lXlb0MYvTE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2768)
K6Wf5t+BGX0XoUvFe6fuLkBTd4dnkkjnFCc3l/jjG301TVMATuw0euwQNbqZh85x
nuHL7/ej2YQDiMvXEBTryjw+1g5X/2G2EwJ33ZtF64Aq5eO4Y9p3XdSRb4PXhYPA
CPBTMR0VHNxq7Qjx0hYLeEwXv2sZStI0muUUReShpLxdBK5uiAVd8soZMfAkSsGr
QwqxevNIVuiN7Ck8+90uqv7ywSPbO+7szjOeaZvzBF11SgPWxblgYHlBrSHjrdrj
mfKDf4/0ll3Eo+02EpNUbKPJYP5vayOpvNotqVjfVmmY0LcEmAG5zjAS745dbwxl
ed3uxYO+NkqYYbe6tyH3/Qh+KTeysAoV7td/hFaDroIzEe9yPUE7ZsSUKepbE/D4
ODHFqXwLLcf+RcXK0G+8btuBQ8CIiGTrpxEM8tCmGFiVKaOkNjq5Ia+nCJ+tYabX
cAI8Muebml52IKlTts7CJH8Mv0GvuM/wR/ayQrLRAqR9h4R9K8slsJpidZvj2FBp
2erNddAIHVbfQEs18sI+7AOF9as+AVjR1y50B9bJnDXqjG0bziNKgZLfOQqQM3HD
CaF9wsSXw7+1Xk1m2ltMSrJwNbtD/lLRouJ5aK8avJaafr62vzTmOBHOdqV9xO8I
isU5ow4Dc1S/f7d41ZEqPfTlDSY3+nswjTyW7DmDLL06F4xsXAA1Ds/9LVp35/8I
eVst9RbuBvFbw0SElyanGQFeIW9fUQZhaWGy95NN1nWfjl7bgX9jy2Ab2HJ1BrB4
JaeyJfPcr+R5XYjpQSuvQhLaLCpQJyUwdGIZqzq426P1R8TThf5AOfisf8R29cYd
EQLFHLcvsPfZmlhwbUQNc2x+Pw6HB0rjdtsVsz5SSMy9zj/bQJQv8g6Useo8Hokg
+gNzYgMBQPFnULZTuY2+4dqwRvhKamWbzKBfjNStJ76m5qE4qKIaP2gja1FIav47
yDPMtPZYFE1MaJeGZyzoKSCvkIKCMhuvVmfrM17boq/78F0mOohIEj2352U35itx
yQVbn98xa+uIV0E2+T/j+4F6zip3gBysZj13UICh++7vMhJi4R5j5WFX5EFIsD+H
OA1M3B/Zgk2k5Tu295oeHLiLK6QDUhOtWILifKfA1t8sslrH7mArwSPyQwO0jAr3
eR+Lqv52Ur+1+/cE9MMieoxN4fSqmUiP6KAYXDNPzmjNJF6AEQv5FcKnbCFhsjvG
j9E1ae5lbbru9VBX1Ri22Jbd9q/L1casxH3KDc/9qChp0dqrrB9+1R1RnBBQcrb1
I8W8wjCB/WcQ6VixJ5FDJiacSOPfcJ4P4YAIGe9nb7CQjQRhzmZnk1O+VR49YDey
zpWQGexD95RDfSjqETNV9BH4siTSHr3fFFqNRTjuViLTLhQeneRgPM9YCl3orNPP
uUatKk5NUAb+XHNRbbI0Uf8N2Zc/2VrYqe+S0Ive05TzEShLie3D6ixeP7+ywctV
65IYgXCgSyIayS4OK0OM0vs56ArXIwPAowRJej5YgXXO8d6M08erWn1w/Oc0ozKC
CPG0SY8fXuPebbx4yPHVl+xBL9vTL65nW2x1QH8OdsUmMChoB6VWBL2bDgu8LL2A
ybKqPwuEweiIML8QKsiLNT5UVjp+quuFTqRQZ4bNO8sT3lbdCT3X2ykaPe1QTt4E
lNIL/qL8EmDYw+uBk40mUhJy5GXwIaUg3/OYUFqi9H66tvCwouvB7ZlI1GC6q77M
9kQHP3c1ozSNp+nG1zvNy7JtlZvJMFIWe2nDOgsF89v94vZgTKU8SjsHEaarHpzt
6Gbio8kiiLd0gNNk4np31l3J6Dt+TJSd3EA+vrMQb+m5n8U2TH6UE79JEyBP4ea8
NHcZbgB0CakBuTfncCi4FyGJcQWu9rC+3fvQupu1XVVLeBZc9dPLRjfnc+837/gO
uQ9d6N95XAQmmLkW9siwI2UA29gfjeY260gKloMGVVusE0/AtPAN01BS6q0HvHc1
6df8onRkhSUG70v8QIjLjFskctoMiZ40gPiZ31SqW7DvuWyH3Qc98fvIxImEnPkv
a88bbTF4XHxYK2aOW5vrLVjend7tbMYsb+tfex7jciL5cRXgdea3vhKr6uLv281l
suQHm1GBbVn2aIli8BG1U092Qd7kw3uO+DspH4m9Mr83Nr0eKHVcsetGKULAP1kN
+zklzmoSEFixqaDTAbeFooUnrYuTY5hf1JPMS7LbWooexoz5f0C8PeucWqnTNinp
Sv4v5s2Hfbn2in1ZjshaBrTXFNrl1QigicMV6WVTzsII9RLhCufJftrftkNHSukW
Bbd90LTZia5UpwFbcgSZBsNoS4ETzas6oXIAQnE7FabFkHbL3Hx4GmxsuLcmcLtu
4V/khhS6dd0dCWiwbMsOF0Xv+svdxNW1YQZ22k+Xu3BkEVFZiCSVxFVvelOzd2ko
T5IEdztphen2C6JdWJZBQ11FYarCFOCb2EpaPFHDZnBUmhyIx9tBC99NsbxYHzND
84BWKNYwgX0YJPK10T8qv1J0538ZBQ8H6R/RLqMxdvS+3txljhOGHMs4JO/3a7Ij
sbixHqrZ8I1Sto1uLf8KKPa7mCTwtmmQWnA3cZQGjceH3/6JQTphxU97YFMglS9m
v06jpRV3N2/q5AyONTwune8PsT4y8cB/0UB5n7+nv820F1QGbc/LGbtYmCDPaqhy
J6VUezXqRHC4M/owQW1xf9O6meWjkDW9Yd6hTcdd+nuQSZh+u6QypRP7x95iRB44
ObKDYqdnDxcNzdIlDvIYM0hXv9dojWxGE2w3UYJRiGJCCmmBK8vKd4O/bqzdEfLW
/5X5BZDLFXncuGxWgLh1PedkHBYRTQGEV6BDDv54PRuuT9eRg1oVnZ0NxB/rJLd6
OA6+tTAWfL5e2Sl5GNQLoa5SzMWTP9FNc0oODYRMqz4orvWL0s3pBSXSitH7e9nc
57GUDVHN7/uRHpLQ7La5wG4M20AP5LdXk5moQ4oHKw+M0kK/nW3hmQkR5QtKtDJU
bJ7l8WV08O3CD/PgqYzIG7QoUNAGXBvMt6zjQQ80rlcYlAltojnWC2o/iV0OvkoT
THY9NV3Dye1zCxCczEEqumAUp8h9Sx5kPr4LhcM88ph9pfIQ+6hm4n16IyRL3xxf
LYq02Q3XgmZhllvwcXHAb1zFh3q3LNHTWJjv6TgKF5Q4dJ8V4bhFkESJ+4WvGPga
GfuR+8LjzO56PLGvYOV6/8c6sbNpVsiOr2GiZ+9/RMjLH7KfHw53WTUbQKq/nHlP
YicrtdrpEOv3ukWJWrneW0eBMiaTcZz7J7VDQXkPWNt/3iPLT232QK+RFjvJD14+
tffdwzb0Cj97tk81Tj4cWdh5wXGbFk/tOqs9+ouutdRTvQDyqw4Zb31NhXngHtu5
yqwYIiIVZYWp3U9CkZCE6dCmomR0xKI12cSznFEv8mRbWycN/2VDrnMU7uvX2Iwl
jg6NonhbAN5c/iYj1UzJ8R6w5iSQXcm9uPCr4SdW9HJHtHv6QZyeZapLWfodrBho
BSJXWGT7icnNR84eBgVO1G/evDG7mLs1mhkJ+L94cU61nqbl5LB/Zvi+SatsTrSM
MRsKtWWLnLThnOB3e0Xc5wGbP53dmWNs48kZ1xYqA4EVdBj35zspmuRVmIp5RRL/
SFwoFs5Vn96zVzIqGjT5PiqQzMwRfrhGa54Uxiu7+L8=
`pragma protect end_protected
