// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:33 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z+jX2EFxnHuOdo7xtiPLhB/i7OrfjGc5JZ/7xcCbPZjok2RhHiCzMbYofvs5Y9sh
yrTvJc9ozYihj9KNIVcc9vFCiwgOMu74bAp6brAgSeLHiM/+qm4RrLBCrdKaNIs3
45eBV8sbvx21k3THwT62swPkC4Rz2DcB0pGdevP45LM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9200)
/UDQT38w1sSSdA9xLEVJ+cKpgAAZB9MmDeJnfasolKF2iM9lHaeS+XvVfuB7eo+3
tVe99J1+xlP6P3VqYR4riudJgYYPMKA/0N+hKF+UhzF++foqASJnwnKPuvdo8wXw
jUgK6aHCKrvH6dU/1On0I3s7HgL3H4O1RziLw+uTe0aBoTZFwYSAZ8vgsUwoVNZq
pTHivT2OpDsMXYDy8ldDrp7RMgp/VvZ99XvJggr2GFlsbVrPfJT+hu11dx38ofHL
q7F5+oYpI2cLzP9ey3gEGOGXbR5a134paCBqqQQlY79RsrYY4cicwEX8qsjNGQlQ
tQQS3mEYRfYihmrvT5LUYtjXsfsajDpPmHkt/fvOoalsI1+PvLLuyWJlbe49lhJJ
ttO3k1jMb5lxVIuNRz/6YQ0f/a2q91I5uYyaCMRZjaK2eVCtTM6JcBrZN5jT9mFl
PsTvKGUGBY/EKqC89MeP6p0OZ8cP5LUsJJ3I992be4GQQnOMM26DH2GQCaSA3Tls
phAaxrVuxAj9r4Y8ItEjcxgghXqe9tfBBrTrlQCRvo/r+Y4AZROAfq/krJiya27r
zAo6l5n6zgnMyUpj5o3/K1rBTjuN5UDx8umIrSpmecPA54UCxvNt5BKgfWAPKWbZ
0GDhJNSp0sCpwPbO5l7mIx9MsAKtJahB1ktxVmX/WWU9wgW9IctLhWRCrlyTrF+t
YpFZVXV1RyGrKDDDraG85QFf1eP6eTZ354VamqRcgYDF3VCiBJLw6D3Tfk44ACGu
r27oZOWVFwz7YCPcs7RXFY0UYmZfIVJqFkeiXcX7l0ypPac8ycz8Xl7435WmhJxW
AuVT6zU+jznCVE3RzkUTphFvEuz7Y78f2x+ZRvQGyXOyv10r+5j9mQxNuC79jQrq
fr2AQxeOYfETgd6DvgjZjf0LG8ikbAimLRw4B8l4VAAit2oyCH9+1d5d+wiGuu2z
j/niln4Q2LuW3qilECce99V35SYs22vo0Pm9kOALwo8Yk8JWL5MwV6uDvEew8dh9
o2dS2ullHOkYjZWLpyc4hfPeTrhC3a5Cjp+aQNh0brr9C+7U1/LHhgxUcIzGIgKk
0MulsDKKooVhSAS29tEYicwO31xEPjX9d8YTdFw4Fpu1LWKvDynB6sapMdbRZfxs
/KO3Pm+HwezIP6LEwyMBnVUd9L1iSs1T9zpPtvgVSWGJ78e2+43+SEl1XmXQgfQj
CePT1uyoE1rZGM7xufomKGJF8u0LaQgUB5PmTFbvgKxq4zblywlH42FY9XsSqnIW
7UeMfFVr3I/4h8pTu87hs0KlXXv3wOhLCIV6FmrvylsDrRfIvE41/On06wyv+B3n
8rsotyi+lxEJXr4T+e8qJcazvK2YVIKXrkzndZsFVOpavGO3GfTADSrDITmSLNOI
G+RcV3BzvMEE0bGk4fEjiAk5NelENiWHDGLyZe+mqCLEXoloWKunLApm7+YZGUwA
6h+AYRuXWWEqsTdpCiCnhoOcX2UFdazbH1eLDBavcCjIpTvyEyPydHrT1z+zBCZF
ayN9nswj/LfQ4pyiEAom+vGjNydRPeUZHOzyfo12G+YF87MvRIrNYpSYRCeRDNny
YQ13wn/QNyr1QFSapDdBzOxHmys23igall1pnyYvFhhS7KSHm36CmAkIUHDFKRNn
cE6n61qbDnCZqEbMiHxwktWLQHoKvmMwuWadO+Iamb96vMBJT1IzMS/RGDy+elln
GKc2jekpBEG4SkN5z4yk4Ip69MwQ7T+4J40YPwKEX/xDOd2nFKQJlnbl2dqI26d+
ae5qiuCYN1+elyXpYphLoxnUO2WJ661CDH3tOsJOshVTYTnR5nC+wjUlIjxfTkGb
wv3J+HAtlaFnv/fWt8Dbzr5lx0urUYnIDEOxk8qfr5lDqHcF2HdVHEQw72CFzXzP
j0KWJzCxHLCjeiwThb3PuvcAzd1GBrhaEz/l/3dLi7DfhFDMLSw4TeLvStvH9Z/Y
Y3TpDRhJ+VnwTQOpnOtK7/7Wmjz8OYvMXYV4avRJzFaxA7dxluUAYAVcYZeq509l
SgADqFNHiEuCUuJEqK72ORzA30AByU+RavgGsAKXELBwVEAesXBZ33XASa2140G1
OqTWarUgYX0rdCUB7DwE3YdavxQAhPKxAYa8D9tOwONga398ySh1H4Pjr8H5UbJW
WAUfWfSw6mIZZJK8pIgSMDOoZ7YGxybTIO+ZEreRGkmRyvqH8bQsK618sq0LdWXS
RVQVgjLnq/7sRL+NTSU20D4Mc4AdnKVmkVZxHGDhEpgZkasHkUqxmv3i7b0u8d66
q+DwBV9J8/lYRHL7oHdQXEc8QMdxKE9q4ihb/97X9Qzb+IVivM3t8E0uXxQ7/Edx
HuUTe+Kp1Oh+6ensrmjqyxJIRTJwaj/+0pcfNSt+0IwkcWJnkYs57ftO9ydqgWYE
gxHbFDz1VmJBRuf33Ta6NG1tDUSB28BVpCcl3Yq1mX2+V860Qfa8cy63Tlw9e2yi
Z/EzekmFBSgFx0IICscklk1aUzg3xRSggPC/qK1deCqbFHl3XLIhwEjpUKLN+EHo
veLtwJNRIp/rG3P4pAG9i4hBPldKZjxRhJpFVAJPIZohePLh1JPeAY8kWqVh6F3D
FvPIF5NjWUElox4y0wOvEg5JY2F198pbjU35Ghah/k7FXYClHEcxw4ZJD4hPerQL
jhaCBoUQuybA1BEYQ3LlhkMYva5Imhl3Y7Ou361wLVXKrjBrsEmXsdFCiqXjLlB5
wf7sOwt+vuQpcIp7+5DdmYoJ6BL6OZRUBTiy+R3a5LKHTaogjSicNlBFIwKyDdjS
lIUgNLDIaNfIsa7QrNn3mRDKFIcVCgmLnWAaP973xP5uvHvC5flPvRGoS2oDw/N4
E5t/bzqx7jjHf9in63bD9qvkCQtb51lzpgSYBSd8wvHRMjQWLx3Vz5od5yU7cuOW
pqbVkru6Nj6gRqO/Uyli72zkK6VLKO26lZ83Td1d8u30jmqVD/v6UkslMC/0MObc
G1JR/ZYRKRBWh4R8QsyO9TTtdNbbORSgq4W4Ou8ML87MUfu8zX70HTjBj9ODS2Sp
mfkgWhp/WgYG4jFNKk9ZIlJh/wyZVn3/3SC18zjnDg8oFxZW1KX2S7C14MjDWmPm
gX4jB9OK0OyNHREI5T8jUb/2SDBVMhrDsAOUDHEYHuqecm0KFWkDSPKZU1vWwzUg
1orlak/9uH0KO6KZ/2SxiEcbozTk8qCJF6l8v95aGhPQgBIba4fvm11kYO8pgtXx
8h3dX2TPPI9oK/fLZeEtKFdx87nihSK8s0XquqQ44FwOjWBRLvHzH2bIgoNI7V1d
vf87d80B5O9vymKSFbXbJ6anGbJUBjca9GHLodYsrFJUA6XKKaZm6gPQm4t9H1Sh
SZY+eJVnEyqTlYtYo/mIZuFAffwPICudk7zxegLETxau6I+3WvWoQhvzMPhh/yDa
iw7vPRcxxVNMWmozrVZY/eqnLNZceaWOXgMIMvJ6Xh64e7lsaV4rQfugvSwXkHji
NaFBZnA39ZpZzJ6p28eXxEaqe0PzpS74MX91VDU0YHwVnZk+H1g+b0leXkXLWSgY
IxGuz/z80J9NrVzfcWK+xoqnhxwPiQRKpyYwrC6HLpPwAdTo5f3jAmqCTQqRnLHC
rc8VtdhqQxGj59T5vSOh8EmK8HVvmfKAMbTK/Pyl6a0WyWrQIXEA4RdQ/EiZDKQY
bxXLB5Ln5UpUE8FgilZnbAaXyyrfu3p8wfiUUJz9UTUO3wi1AHzomlJMVDEwp+XK
INqiCTnaTbKzEq5Y0c5Huk5oDG1g4oqeZ4CHeyHCu9b7gkQJp4cXyBGiy2B8SLwC
J1GN86tTPeWv8kjGc3RM5wjCda5YGLAe8FY4E+6UO9vr14kGd9ab05XdN5W6aMfa
HAZKdcZJEll3+dXag3a2S8DTEWcMqCuiTvSw0Wwt/nKFObDZrVRd4XkelgBBgMto
DEGiPJWTg3YpgIgEA/m78jScFTDFqIlO1C4RVHVzQ6lbp6ntQGFRfERPLSpf57zC
3MPbFoSR0UEKwYxSgnKCKXshE7c3mjPAsaX9N3L/eD9pHbUcxmVhut8bxnGwweqz
JPI8So1tV2XBBgIDoi9vItroWTQn8tgjW6a1/namoW/zKLpJKRS3Z2Sszctz5l54
WdpZM9eyWYSZhfzdnZFHyxk9BRk/r8AZpUvZQFlZl/UyBVEG1XAmcBLsW8lQEKKq
1wqV/qCev3EYM6gPZj09zAqcqtDMsDI+Pq1miaRrSuPXlEY3hRw/SBgQEAUEvXim
BPzBRsojHPL4ILUCDca75WwSi/e/nJqKncIgDW05OFQrN0eQ3zIwTe3MyhkOE4bX
s6maOxSO7k1shyhzEsyiH3hsjeIvY3tkQqI05tn5i4W9xYaEa2MAOvnr+6Qb+eGk
/3sb+vmQCwgBtM/8+fm5dvvyYCuCnng6Hsxhh+x7rybizPs+kM5ovKlXWQaTdO/X
lKNwV2J4FnZ7+JtlA5j9z0r6PBR6f01g5oWbpTEJJvJxWVYkP2OWgwswEHyK8gpq
W7C0R1xdPKpmqPSbkoVmdgKs9HQ7tQP6k9NBouk5rvsMxbTfEGGESTL/hqVoCPDb
cKoTP/Z2aZNTRIDtGdw6eohnHFfw7ijMd4ZJxg0I9HIE2FpnIZkwEZCJEZXAA3F9
TXliYm8buMRfxS5seL8Ek4AwqD8bNo+7v6lpwG9yBhmZ063vYQbDmvbaFT2MMG0d
QbWpJcCn7QZUdurNNTnlz1CjzvLIyaoyp7SLxmJogIfMa/13arxH/an8Gs+9Le1a
l14/Dfl6z8bYt/VpF/vEa4y5qsuE40LBTpv07NCRGE3dzEkajGYUSAoPK11CgcTs
mewNwmcl6C1xmWiYKdmezqojdXeJ5WKB56Sch5C58SfL/PB1/Zr47shGSRHqATqk
pFJizx6KRQxvoj/H+PmF0nnAtYZLaBgay8axXc6G0DVgfU8yr0dyIq8W/gniFOpJ
k9JIhQcADic3DthCbfTrDGnoEUoQP0h9Qq5xfmnjGvKUozwAG1ntBa2fXgZ24J2/
UPgouxXUwydhTbZAp5/th5/8jXLNWUclTohFGwA2mbXLbRbOC7qsKY51WJCm2YR2
tV7aJVdGCVsSWFO/xBni+5wZeQgHYeeBvMldlLbsEbe2otBV99nRpDuzzSGQIAKt
HQVh7SNiwNkuuOw6i/mF53ku+JbJarGliQOulPCyfmiUw4VdT7eEV04BF4RN2Aox
xxvg6bn8kVSmIQ0RrJYE2GDu72J3PRPFSNaZnY2VvvhyjbDYhQf0J02ym6vw0UZS
3wac2SgUZ9UvieMjTPV7Nl9ONQ5DHMt4BlXtNqSnUP1OJTl5MOhRR57HTkzW5QUs
NgJcZ37pOvsYWu5B+73Tc/weiLL3eJP2dpFsYnywt41xTucUjCD3Ix0/aNqXMenQ
RNOg6E4k7IvDTkkTwTOnj4bnRmOxH9qUCR/CpY8DZ0tT8l03bxSmdCpv7hmKthiS
e0CCGj14cUJNn/XEl4X4sBrtCa/ppNB2FZxqHZOTip31t3dQ5N6F9cofqzRNjrxp
+gJXFWMDdr/ua/s16ojGsuWfKnmUGMDfPZCW5NMb4699rbU4UADt0dE9bPF6vscJ
0CMIxcKFmSJr+pPw4tXV4rpuFAI3QrF/oRkNQip4XoAGda45p+3z2HTMfk/4b4QW
YViHjiIe0qFThcPNAFgsa9l+0QsHv584nKHW9C0F1uj/rihSg8K3GYCZEVfR/uwI
uO/HDRTloUApUe+HfykEpKRs3tX+I5cOoFPQ2AHh80eBE0pP8+VIOGPjPn/pWHsT
Y3oDjCgmrUbSzAEbYZMrJUqSIpO+2w6N7E1o8BnOQzO+xRbJkhrk1aYCBTjh1KXL
rKFnipnYGnKjnEf2/dPT+olk2YB8dJjmmapsoOou4O7D7g7gvAV12KDGpRdeJ7kX
fVE7DiQbA299+pzH1MlDAy/5I3OE4NHmj9YqEdWkzdSxL+0T8OZSHCr+F/YauFe2
OoVI1uIrfsZC2d+p8YX0QvqlJfOXECgMF1vyQpKqwm9nDmCkA44PUpPSj0xjZBQS
XQpa8Bjydob3nVQo7sG11IKrUiA41/HqsmjgqFu1tx70CjasSJsAQbUyxD5oV9ao
5QOcodMapo/4ANrLJP2S7aHPTJQenhYVpTd7Db3gexdq92wBKkPIIEINrEh8cKFU
4QxN3LF0K5ouFT6dGmp09XdV2ITxNGebzCRje65YSDEVd06DHu0SyOflW5iN21YE
GQG+BcneSFBIvuwAKZyXt4w6Zh7REWKVHPaQoau0ZgEO2zgiEqbmpKPRb69qW6HC
hTNgFlRAYpA4C464jWTyiBy+2KAxE2d/PZqJXZd0ab4jQY3grVZmMUyu+vcPBonM
36nnjBDfJqzw0Ao+xu9RQgCm++/HX7UJhMYfQk0MTY5rZCQKTdyWRinB0PXQjxQm
zzrcjXO0HvA6GywHWezH8sPMUc0WX9ffgiRf32JIglZVly/4vCf/M0ShEaZCPPU2
IqMZtOlyJWvIqikI5pBDlSjt9aiio+jHbNwUciA0Kar6laNERu2LEmz7U6hiFJjE
nB6m9LSE8e1/fr8JUqAfODUiFjbhkrchy1XvZsgsKV0x6vvUkV3ucua1Zl97boNQ
ff1bPRi90l7NNAGmaFEfAQ1in3ej2w5IzhEE0X2gx4Mk/6c4GGMbMIS94ctd91lj
4sVkWC2TMdFfsYJv6RxQOAYVAVCfl64FSC6zC3fQ5STdieqmakPUEICv5hrdDOlX
3RGkql2Vx9sY+tC5Ihyugz3VF/B6EUhpi1hIKwSTY92tex+x1qBp2c/jNFUkVHG3
OvocVnjvt21m5FwkBW0wK/rSPo+TZ3RqD3EtjsqeNejbUQvwYR2T0HaaPyUKMHdP
Ewo5jcXVeRfBzAfJpEGiTycQLHmqP161Ul3a0TQYeCPoL5R6odOLSumBfvxC/6sW
BUWeql5tyjLuvmwK5Fk5HqLWp46eV7I/pv8jisX5J8qdwJJhnt55eEhO5Gxa697W
64idTbzarltO4l+m7Y/4K++EA5AeUMa7JWSa1s5Xuz8kdDvwybf/F+7Fl4ZudPfX
JS5Y5E38gCm1u09gf2tpIHyfnnYo9lVJVLmie+5ghShtsI9vNmMwUT2IGLeG1/FW
YkU46HwjJ3aw/ujsEEa9qzqti5o/I6xcRCVkc3JgwFswgrV49WibBxGmvOB5AKnl
IvtsomZDxEqW+tW3105qWPULFJc284Ywe/uXY01wuqVODJ/DaDzJfXWABQrGRcl1
H2uurRUDvCvTisPpH5ow3lCgNKONGYNCqDFKIFCGKL3gKeWQ70RwR/ifD+jspZ3R
IOBuDwD7eMDMnImrOGPunzY5WsT1eTsPXfrR7F0Lmy/jpabC56ux0xsWSt+P1ubv
abK9hdvgVX+5+eByC9MDVRUAvJLIvccX860infpTQ/oSrM8dFu5jN003XkCUTx5q
nYIqncC1J7URV55VSj9sLzca3IpmeHiYctpGbSbyN4UmpKaYJ9qfjYQT+EA5FfH1
x+eVlkiP6pAZY0+jo8Pag/CAwkJ2IxQRdvOSeZUhkIdpqcmcCYMAHG4QgYTVliG1
y2yAAUH95kYuxrLbcA7TOBfRBkVJZkb7YYkZMCrLU3PnZOMGRk7KOz8u9/niolGU
JfkYNeCsoBkkXnI6RPjLBjRWJ2OMAw2HwqApLml8MGHyPMVmcymX4Hfgaq9nepBD
pDT15hk8OLQq4tAXqsEk3xW87IB7rHbSW2UIuXwqUpkM4hQxXmodPlqhvp3BONnH
TUStYb79kv9mDnvmcQRkqa0YHw72CbPztsPOi1GJGPkZxfZn1ejokXIWXaHVVRHQ
nk7jeb8jNdc6Ve5RtzKSDaxdSp+6UifnZ5muJokS5Wem9sUDq/NYWBcZ0XfgczGM
2q2JJJvEPhZYLmqv3zqoey5i/YhLhKov3Dr5koMVOknZtX7Qr0bwpOcPgQfrX+SZ
6TYK4aZK5GCrMAXGidh35tmFJaxv9BKDyg3e43BNFHdQDC3K3gPVEeImx0IXg2Ts
xWBbwtGQ7I6wVA7bWRbe03V0JbNb/ybfwBydKFuKXWC0u728vqEG5G4lg9mQ2kpz
QUPGW43GpIlXBdE6UI86/freBoEdgzLF5Ay5J+yiq2VAW80sC7gZlfrllFxH5Ug4
PBDKA1S0usNTNHByyDo/Ikcrv1nrLFbLxbJoSeHrJ8YkW9fgAjtw7jrRcTnoDDJw
U3/nrzySZ8WsJZnRcuVEY8HUVs+lQGbcAdbSD+98aaezFYFDF2kIp8NvFzQ1IR3U
yRyapQf2ImSGQEitfnP9xVItdPGHxefxYGYVfSvLAe2szFASWgTaJrVj484bIsoc
7Ik7dY/CSPdf6zerXrWxhv9R4WBlgGtcoSZQgxlpBAJJFigO98K7htiO9hp/v8aP
8AIGW/Wnz3cXpYGURst2xlNZi56G6+iNEDNwClZiVMirywvw9+pYSb2TkQyzOCL0
gzgoCO9eND2Yq3vdqRpulsj2gQ+FFOlfjJAR10WcANzy5Up6WdOag4yY99HYVqg2
Cgnh8cAnVprptsuSKmEuk7fTBV+cmeM3iOqOXpb/+FzB9BA/7PrXKv3Oa9VUawow
FTQxYZivcFubqvQ6dI6e0SLVMFb7k0X3JghcPYoAQZvuLJ9YEflK5GOei5c8zKU+
EJbGi+8/u97MQIRvUfUe1fDbyHhGg2kN7/SwyBTQxRIt0KVR5s9mLy581CUI2uL1
KUbqZ5vniw6Pdssi1TrGBFbiAhGK25ZCo/wEvqyhDY0UBfiPHAZr0knvCJczPn8v
6w4pHkXYdafLwB1ZhYjXwzFGF72Tkfg1MZcAqW75I1HSCct+QP6QnfvARTd2kgIb
8QbV0r+dS4a2b8Fc71eyigJ/4Xe1JHNmwnuHaUzA07wsOJMX1Y9px2l690w2lxT4
6iLkYCbVKQLv8fZyVkHTTG7BY5DDbeg+mifd09T6F59c+idFquNvOJtB7ZizOJWQ
aDazOjv5ViVf+Ll9bc7E3gJkNCRHae1hppkrDUe2tq4CVqnyb4vnhDz5ivERhaJc
SQoif6t8QIt0P/Ee1HE7+/m6C7Cdar4HF0iJawrKPsMRmq2wmU8fZa3FlIw6M8r5
fqlDeVTpSmNJXH1OmIUmd1GAM5h3SJ/GuhlQ5L8j6UBrJ7ly13YiJDtdlSeuEYGc
CqWTfGI3HeXu5AURhdyQ+ON5UtHMDWfbH3jD70tjQ38LEGgfppemzDT2Kr2iULZm
GggdEFWm6j8MFu20MNkjmQv7lrllbHLa6qgmJrjZF4bovkpbVRqdync8n7VpfpgI
cYG8V8DU3MvcNNy7dh/6+bmEDM7rJdSMyLuI0ertR4IeSv2zzOAhjszFTw1no7f6
/qrGvbkTNXBo/QopyyNltT7tYm3Su5TgLhorW2dzQE90YI+i5pkkJp5xXVJNyVpM
2XihB7CXJrVWjTxQxa4keazUgGw+/A37tITUpENIxtvPIjtLXmzb9Um0MvkaEDN1
xA02ctsUlWgVgNtznpqkmO+bz2ynSGO60QzYOohmhOxOb6mddQrxc/W3yl0llbmc
JsL9xmmclMjR5CfbbQ/goGxI/lo6t2HRqhKASTe9Wn/+e9MYx/DcEGZLSR/jhqRH
X6zvEbftqFQ58sDicRR3XeJpcPV++VNhu4kx+QBPaJ9LXKam300THrU5uuoR/bH3
zm6ZB7ibik0a6grngYSQ2uwQnwR312TS4MnGHGoAxE+PGL5ov3zBbVDm4GZFuomX
4EWkPalD59+mW54MeATTRj1aal7tnDRMunUrTAtS5D0mwdCv82Xvx3iGZOC4Uqx3
vjG74VhXAtji6wvp8FYWYJgMj7t+MtStLfsu2GYV4pXrgNGm6utRhzmttzTW8PRY
B/+IeJmcVh0fyDGxGE1eMtPKH2jVDUk+iXZBvF6XyVsvMTWjHtEG70oavJJY6FiX
FfZxga5pvcmSBSC29AlpvQamCgrQB6reoM7+fTpsWegKJDD2zZWvntF6WXFMNKSM
vykt+q13ZGoctsiqvycnfxHOxJHaFjiDZHrxRIVK8vjrIOxUcvtJhHfLex6phuB8
Mbn+M7pCvW+3TLpN92lcRDjJQxFCJV1arr9OPab8NOGG7Pt5ObeipfADwXo+IMbQ
9wBvLs50C4itkbflCIQ2bpjnJAfYvdYlZfjSl4GXcRHPAith6a/rm83gSTZnrVb0
QQVypsbBJTb4TGBwPxFudwchzfvjHzvr+XAY15dpG1zklcsh8ld9OXwqd5Pp4ugW
joOZWMsowCxSsM4hg+H8t25hbfOw/FZbDBmKddTO9oWJ2b5qVRS/ujgGo+6QRiEp
PgM3UH0ekr44C8YG8x07L/nbrlnpI+EyTMYzHoM3Wa+JbOoRnCy8WJ7aiXNRYS/t
u/wXR4DfUVPQpSx3KdbQb+2mm1I9yTEMAfLhBcuyEFCe7JEymWAsPe4VMSfA36Th
oNUXraUllhjwuXEep2XqLCF7vqe+MmFNFKpH5GBAReC5mnpvnVEnXkK3YCmKkx4D
8ZBh4f7q5e6r8GUyJuimVmITkQUDblWtvywmotEU25K0uBKddRy8u0XWavig+yuQ
9hMR8ecdU2/v6KbEbrz7ToRIgVNtpmnvWn3swUrjFWUM8ClP+uCUN/j4Q1JF29q9
+ICT3oJAhXa4jZNE/doKwKAaOuyubolrDEUUrPajJufwTxdh9sRH6FlqkeFFLPqj
z9i5z1q4adk3/Wxgz8WKZDCf8ZR44hnj/0pnyN2aMFStNAJfiHKRd/q9O/WuU978
VlTUSuCjJ3ogGkZY2E8/ocYqoNJuPr3UmUCmG6TQzPxcTdM2rc92B8o6Xcj9Pmpf
niKbFNXNfaKybo/wghaO4mJtPOhoh+mEFU5s6+9g7ySZQrzltuBoLWgGtlHCCXv0
3bXhzy4koHC7ot4v7UL2vW4xBlkE+WDMMvhXbavVkOQAdlkWkWxCMw6eUCDTLuTC
qj/TlFp6SDv/WZysaI+R/buDKz9T03BPHepWjGiJVs9oLQvdcrk5DLAlA6gl5Ncq
tQqangdFv3K2Wb5+wK7OIDuCuUXxp9/ez341sOI/2vIMoZXq34VVZTVw8kue7uEM
a/toL7iWYtCa9MZpRZSM+Z5zoXcFGY5x4hOu7Cyu+0pyLJWccWH7aBhhWrIQNH43
Dufvxlwz63hqt4YYDtAn1ZHLae4dN/DLVbeD43mJG2ffwMTximSJ4lxakoveo3Az
/rKhj1YWd0/9ExTZzy2Qang2vNAQRLMPQn/tIpdbpBpjVqXl6+eJKPxDdjK2cIDz
xz4NKzVX3+f7i8FL8u203kr4EtLu4wtC0rZ4bfjSyA0BIYO6gBsOHRqJI2MPyy+p
A4UpeYY+DBsyFQhYEhwzPC/XThy64+FL2OTUuNDpvkjhWUZWEMRJSiJuAt6saA60
s6xjy5yhaqnet+T2cO/eVQETNap9CFBWyPpY0WSrAWZ4XFzNPyyiIx36vaGe3x+o
f690NyLB7s4fmvOkK9zr17jxDZe2tLPVn1tZ5WDyC+mCwMkyo4y79H/TYogC9n2M
5L1rZOjY2zaSnWmdljxZMB+VpxPoaDZMW37sZcHQTUeWbzYyjZryq3QUTsx6judv
voPBiMEOmNv4rZhZCHDNvb2Xaz2FbvGcWwCpIMXck85XJX/2YwffbAdV8NvTlCZ3
TBOuD4S7Uva6KESaKkFRuC9/qhP+O8xs1JSH8fTn4wt1svfjMZkDod8MARl5wUBz
CPP0Aeb5Sz68E73sv6LGF5jkx7b5It0Zxx92zLDJTlSpWTAG65/gtTJ6zWv7FTS2
4rKsWVaTb3Iw5JwWXF8d5XsCbmSRfsYCbAI7R9TFeY8Gnb6kQa2n07fs+ZRIOA7u
yKQRMBBQmfulgVGu9TODQCEPcrMn3625+eBGASyZrgQclCU1igV85V3HTAU82rsW
rR/3luEiFecfTguvuymZFE9GqE2fuUqFI4jvwA1xdbmUbejWLNHNYXUMez8VYqjb
NjIIg0VtZibfyj9grePYX6f3WVEQY5w4nCeeWV/aD4kGfb5wmuHxNWgLyUTWlt30
N9c5EFWqRDVCOJNsQTEcnIUaad4kKHNO5Tvmhucqd87dP8Ko67SGwLmONL+yyzvf
PaGvuxK5qQxFQ50sdMBoVZZdr9aFCnhW1/tK6+UL/oQTJ3wVdRGtXWxMX0BzJD/z
+2yLLK44skRVi7SikzWaCxARU86cydmcce0P1UY1tGc=
`pragma protect end_protected
