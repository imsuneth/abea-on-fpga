// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:45 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YYYlN7JTKoFZArcPyXLoE4bxRYAZQh1mrORGZBmlGxz7fkhyjnjkymZFNuZIW2mH
xzTIE4cPue7WGwZz6sx2vGIV4r2hKG3bKoj9XYHp2EwkTrLzNGHxi0GZRaxzJLS7
VHnL1BDx68VY+XwZVk3mT5tnZQNy38qAxInP0EF2VnI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6560)
O4H3TvAjjQU/JXCg86yhMHMGtqvNReo/8Da93bvIZAWPMSWSXHuC1rOJpjR1LUrN
W40WPcwvizCzeH2ZsbwurVydOeZ09EnPz0VJynGzjX8dtnz7z5immUE0HNKdAB67
AV4F2FoCaFtPvkjxoL4EicOquMcHjl1Z3Rv5wU1qPMVFO2ixAlJJ0bDxkGDvh4sa
SIm5Mi0dmlvl078R2pgVtyR6Q9pXC8Y0+4+PzyoU3FvrTXTARi7KXWavlnUTl27Y
XWd+uNup43tmoS0pwLHesVPWPWFD+um9FCwIqejeosDNN8PLZxd2E6rtlr3kNF8F
PuWnJ1MkjT11vsBazURbk65crL44wVAvIUac3lR+f70y7mFNJuZnAOjpPjsBPRNC
c3Jn/jFe+5R5uNdT76gm2qlqtQacvKPHsDY+UOQBgOyrbWrgjG99yYSBYJTuphBm
5UzQEwfqk5mDiNsioyKxzbT/35GfaSThL4x3f14xc6oDyCFHBuibkQ8EGWgqnR0d
L6vT/xkE0+vC0XxsHc5ds0ki01XWimwpozeyU9Bfm89CtaMjbPnAIAe/p817Ww/m
+4T3l3R71cEjLkbH3QWSaxyrW4RoVe/tHX/NYmx19oh2FpQTNkwV9eV9ArD/6k06
ZZdgmYl/CV12hYa5kNi4eosRcp1s8ijFsgaIhWK+jq9+MXLHblEcTx6njPZSQ+1W
WwcScZHsmjHzwpNdlgb/0zC+cJGF657hZ4FUxf943WxkkYSL49ffxTUk4v5KNtXA
QLV1TTGB/+sRXi7+cn/wSSieNz9fM2B3U0ioJ5fcdGpK49sa+VvsMcR6fXEUyQZ+
6C6GIqqMY/V+8Qeibd9SLBL5HbzF03ogU6DKVwyaoAvgx01q10ZTAvWVk7JfvfPt
f2Sb5LXP05kjXMIhjVqQQnzISuNPSk3KKb+B6GYWsH185J2PytaLg1BSwsXDjcTX
PIUIs9qaNoBYn/M3uPyddkPUJkGHKIDNqvuabGw6nJImv4NFGzn0sxI/N2QvDdpt
XDD3PIO8vKb0XhKLBpuTW4cp5c/J0iexS1OsIXjgfvH0xMQREIZK1WGU2zgpA1Et
b30nSPW0aldnqnja0o5gLa1Kni9coosGzL/K0sYZ7AVLg9rJFaQKiTdb1aDt2XSk
rIlRsd4Fw8zHWi/BSAkzXCWndMhZod+FmqF4LVo+qxlhKdo/tiLmZixyUFUrgJ+N
WLEwV38k3RiFn7arGhXFOKEAsKtkcmfyZID4XEj3NuzbiY+3nDD1xnAQWT7SP7k/
vij6gv8+dagM0nC34SkCGnGvYX0b3p1Ml3/rhsVFR61OZFVR8BaZjmU1WsS9roQ3
2HlNJ/rOfC40l4Bs+VKC3Dx3n1l0murntPq9cgs56fOUGg2xyOlsk1Envh0d11Gj
TKERUT2Ijv6BIAQl5fxQl6xLCsGh+zvgDdLri4ywbnz+Q7UkQAkmZKAu2SkY64Lk
O6KQC+t9tJQA2h6NJgitHYm7wJYBnRUiydwTOPmBYgAgCU5aZzVXfYUIFtE+Y9lo
OBsnRIuYgQuvxaSGjUXVifWdDjkDZIsqduqvvSp82wtbuM2e4vXpobvQPNiBqvyp
U1CG6Eyi6lezE3oiobcYJhJgQK7fZGjyeb5xdHDZJXLc9hKGsSr1ialR033Mlz6R
/wUP7j67p502b8uCkU+ipPHrOI3oLX/ou6eH3WSPLB/0CUiE2m4ez0KV2A7Z53XF
T2AGN5JTvxiTJKVCrspUFOf6L+NNNIw8LWwiDTl+XcjQG14oXsS7dNbCd7tPdBNl
P7rX3Wx3ug2aZ1gJ4lcmGl78re6ifAJCnT+QiBChgWVYray/cNOy/rVZ+wO+Fug6
/AawP90Sn8J1Hv3UXLooLDVcojdSbA86muMbv5vJuQ/snja7lLtkyQyogkoYQFiq
/Mk767oWzYq1qelDlQlrysz9jHdUJl6nNXIZ1T/1/N1x+Pa+WCw25pqsJDqTXAzo
AGh9OdivBFj1jIbmOgJJpBAqce5gRUT20jMUriOCo7sZFfnvofDWmS8fjwcUoIRL
0bldOe7mhHIXJPDWVr5MAdAefncGgGWjEmOF9o0eRor+iseOPkrS9LnPESqVS8wb
jI6h6yVgLR4l/7fqdDTL8wJT0B/XxYXfwbmBTTZQAAc5yinnkcHwCT6CEEDYFG3l
8tm9fJzyo/Zu8XOBu6fAIOkR0Jw3bncpZJxeIf4qLFHXZFJMFK062MUgWDxsgBwT
aqjTvvwkktuIhY95+sBLRV8eFRyDh3Il8x9J6bXn9/3hnoWfQG2uHf6lMjJkT+DC
CdcjaPCKPAe/7lDtCiqNN2tgmeha13L4/mX/zVxMLpObh1ob+2sGOE16z0vzR2zR
AOcMg8Yj/VxUBjY0I6rDqtHwLUjAM3QiK8VGfZme/aGpZjjyjeZfKHD7bV/1rpGo
Fr8wNKGSNZ0r3j93cdsVg1I297rxGhQjprj60ZdDdf2XUn6RswNNfxE7MJ0MkjLG
g0mgm+3WFjHJY0Q2UzlURr3GtbBPviuGY0Dvl45k5m0XF710y4x+Rqdrg/S8ZnCP
CkAJCVLF+cWuqQaTKQEOkWlbAJ7uJWuuc039j9uSctTDHCBqJFsrKy/QT+vKIN4+
fmEFdbQKPraPK6daYuV33G729A6xpo6xfNs1fWH3a5P2OvXRSm7l74M7hNkaWi6I
Kcy1cT9N8L15un0RoFpPCsOXA9mCSH6br2A3XgxXEZnLbIGZih0iwV9tB2pcQyzZ
D5bEr3dEY2f8pUpYbdv+pvhxLK7eLuGKxsrNtPpsLj8D5DPGItrQYk5k5dZ0djQE
kP6eQ1DkNDYTuKDgvdiEQxGM5lU0BMGbrIYWy3mpLjdDmte0z+w8VewjzQh4jraX
wEnJI8oGbRMuYZFprfC6TOGpjWSIImxdMYrFw6NeJutxk2elRV7io8DT2ARp8iB6
iacYUWo9UBoRhkLP4Y0cLIo7admtYYI49y1zACHquHuyTM8crzBuZDdoukLkHIAA
TYyO3szHZX0coKRK6yxxHzn+Fz/HM6THa9+/dSDxcS2kaek6FtWwYCrqW+AyA7wL
nKBdLCv97wyM307d7SqEgPhyf8rpQmuWEuMcvM4fzEDCwRy20lMkNVqPBCgs5iHl
06Ljn0N4AsjB78PV4QVJPLQWb0PCx/K1wAmZGv2XhKh9KaDFS+WvCE1ijJAuXz7s
CyMsHbrQGa6PecZFuaWn8ed3jKpXhZx/cIpQs+RLn+DKFGAWZTVSgPPQo9Vc3+da
N8TG2WwRR16AJV1EEjDeQ49cI488G8Fe3uprt3AgzddPbA/C7Q0+s/EfTSEmvNLb
tJa7qSYkK8Q4ysHWnWO+6IkA85SuUXPsmSfI7fJrJji/EbFFsbDFB4dH0cQ6aEIf
bkD/D1vAf1bHaswt1O2l9X4Lny/vghFmWWhZxqNwZl7Y034C8fIFfuy/Wo4uGetw
aQTe/d343GvDIibM4+zno7xWF0l51zSgT/KRWmB7mdPqmjGVnYj6BMPbslz4UEqK
TPmTk6vOmdjgDlzDeGurmIDFZdQHSOZdkTS7J2qaDbJC3HCSaKdNgnLqF7nVtKh8
2U627giUIhvDHyz/2mcUkC/ZRdo1ZezQ/jKeZz+R1VYkYQ/uFsdbUhLWXz1S9twe
FRhkYK6HH3dlT0tBJ1K/UShEriy7sFonUlOafONbgYkJgTo/hAiTbciAS7As7/+a
mPKuc8cyLZd6zsEgIKBXcemA+hDfv0cCnGAySfEhWaoreJffXvK+SQhrMXHC9bwr
QD+ca8Jgi73mcsf2RyzPgfk1rSfo68eMtE9cxsKShlleGFhwvM+p9Ttg2o1Wlllx
E87IDfKlRQUGDkfqN4ps06CDoLrNlip1huei1ShAobF7ySmF2CvyN6w2ukfQC0Pz
2WhKl7FGwt5KHI7RZdB8ehkD4WkEa+swysvsVQJpk4QhMnV3eTAyODqwaMIWTKM3
XlAuVLiBgDjF56+vX4rnfRosei3HtL0M9onTMW7bPWV+3/2Y1fd01WNcRepI93f4
ig/I3KFz/gWH6MMWozJOG6LK8bkmQGH4w/cwfnsQ+yQM2AZCNbCfa1OMZYMkQHnT
JuCU2nDNug5TzJamZqSC53RexU8Csm7By6xsR8M4j48b/SjlZT+kU+qR5EwlFqB2
CzUTz/NsyY6USla/uiUwfo9y4m61Or6Ku6IfUAfF9Vckn7OXLDEBBDfpdPuT9Jng
Zsz5wFPyomkKZFi7g9gMLEjhN+w8aw5pyZZjL8gYIYhszwSP2gsEdZG5+cMP/6f0
LR4f4pQsdVlbClvaYXuY59021XNjdSkpJP/67/JnutLneaJsYUA4YUC/i4hqeen8
zXq1u1PCEstGlbKQdvYLhpQuoDSd5O/TTVj1h3fqcWm0zXGPJLGpA+uacGu+8G/i
T/kyWvo7yMqu1Uu9kq0N37B6q7Br+Qudn+Pgy/NtZHqBn5OHqwxw+kwBc9pMjg4k
u45z+Hq6cmpkR0z4e59e6Vx7E28lk8Lj4Zwdk7LOTMUafBQwveJaPlTs9qGCED9X
YzqOXT7wK63Z0tMQnkibO0WAmDaGC1nmCa4TimgIA3R6JGWB5IUIOG4rLSK5axtB
Hlop7/evfYUMS5mQmRZmTLaaGWccnIUvvsiPqsd0nFD2fABqsOszFEiVNGCo8bOJ
FJv/NPzjBgwgebJIyzNWMKW7XSUzWdZHJbvUM9+lBQkQJq59pQdcm0fQUT9Y+PfM
s3CUyNwJzS5jgqrQ9Pn1RTnIFJ9ElSFUNMHUMDYprKFBKVifDTdcsfhxRtIW3pcS
1DRF9gw0wHC8IlOnqbKkIMXPW4mfBZ1ewccQiE/gUVPn+3CVpRMDweNzoefR6cdk
i1N4IBNPK//rOP6vY1LQ6mK3inE/OKbJuRemmIclWrPIb4cmJJmBf/XwmDnETCCh
e8XJIBL+YuynCMqaxy4CjoqnU5NlcVqOIuvlSbfiGIUhmJBOqCk9j/zhorYOfiQZ
wAvG5Iz/3TNiofVq6KQxnqeliYd0lgzbVL4crspR5AcAmD9PwgsqAxM3QbbQe+Jl
bSQU4yVS1fx83euznE73Yb7XVpu2UVAFaC7qwz7n94ne8nVJrUfaI9BP2yOxENWY
9eAmS1yDeaIZbHjK6pw5N/1/T3FEzSn+uHclZ9YiH9n8KDNJ7Uil1oC5uPyCMs0f
e5fXFL0E/OBa5yK+xISqQ/syON1KKVybRf7W60C3b2ayBb3z5FGUyi5XLLrh9LgC
eyIPBRtx83so8teDJ1rvRfWvprir0d+8q+UMggPXInbLC6S73gcifeeoLg/KT8XS
Jrs18hPCzAr8yITaCCk2NrTqCzOZY056xy/WYTAR/fNHK6lzoDTZYeO6CODRi4On
FZZQSX6aUFlEAzbLpAOdB6c7Lfnsxc9fcyGpRq52fxhxNQtKHuNZUv2nBHsEQHn9
GXjKV6HPMeAFHd935Eb+zjWisXK0omJDtmKFE0LYvIjRRJrZllRzoP62ZgNnaduh
9ozwZ5DWkOW0lg015+HMUuv8ud7BQ/XCx7xpWgaiup79x9iXTNaRmHfQLpQ9VNhO
F553gp2kVqjBHqqTfI/3UOmBlu9klB17qs3pzYysgCuxsGW7AU/cAIbaPYGnqm2B
KWCOnML+DoYqFInbIhxhFYCqZNC9vX5KabuIb8OTN2/3gXCwxoM/LClsjOY2aeqm
W1eiDXcTUOmliC1BbKYaDQKqOd2QusMbKtRjsHnL4l/Kok0OPfQPX9ZxqfIwTWGb
NIl5inGO1qp0JX/IK0b/uOQxjgGrfplx9sL6bTVpf0mubkmU52Rzvmbz2t9i0KDw
AX67IxosYlX5mGwS/TyiQyUK5I5KuXxwnuQnrv6xl0+95vXfNffgF3s0Qjz/aaOe
js+IPtDvVTXNq/BtjH1yl2P4RtpNHjlEDC419TBR9F46cve2qdgKqP1KrG/vZeOR
Zd0f79i6H3SmPlV0HP3midrUX7iXHPem0q9TF+JLUK9PrnjH5HxXdlCL5P1EHlxI
fKW4Jew6LdIK42J9DHqq4IdK7kStFGJ2blbMNd3p7RPcOpHZzYiazehfhxwNgaJD
rlRbaMhnRfcUTtpfk32CiDtyW0zLqcz4HSZifx1TSmJLE0kmXOBfm4Fl7ftramwL
2v2ucw4vI9gz9ggbNi7iblk7XdPJ3rlJyOnByEiiqIstlVIpf3TllNNQx8gV/aw8
f8a0h/YZdMauakp6qaw6HOLFdyMfG1Zesw/+MhrMTWX5ezM+zgOFC2jRb6Dg/M4G
8QDr2mWNdkG3hSWisKaOVpE9xRjgTo7H6pdCBFsG8u8sVDjJu6UWxB29mnK5//vk
pfPAb4zXxXk8Mz1GN9QMKj8tvf7wlugcqlj52Xe/77VZVPaHE/zo8VrINLuOTrLE
3AS1LL6Yxwdf+F9UnM7b0jG0WOyQJeB2+BajOBeFM6LN0ZjimbAPsQO+k3+k3dIR
t9ZNsmzw7Nh0lnj5D/b5LqM2vyJme+iVaB7tIK6POepBSwzx/O/x0nrSECsISrw8
oKaoXI6zHJ861wTylblKe/SBeSNK8PFf6BKfFz1ruafcE2k7eddQetU+9Fwqp3gx
mHLC3pXeLnGdixfGKHFySR/XY1/sTbixbc3x+IDUIBGT7IVZaEnoKrZsXu1Wf/Mc
pwh47+/xa4vHeYiMmdUv9fB8nLFscXidIAlGbL6r1b8X1j3K/fesJMs81Hi5HtZ+
Et5tlqUcegxwzCtxeJOt40+uIC+/6HI9BbOHQ6TWkZuimQLoSa6CLv2espI01daM
rzvLfg8xA9RUStJIqvwkj07OeIxfgEOMJ2q7WD3e6VqCWCK8faFWTyoZA2tDvBAe
xoMPO79GVMq0QjHnCS8omacIPA7ZoWcCI+1Hwuq1pq5D38qCUHwBcW+UD2ibyxT7
sObvGkGx02hs7gvSatoYarC6UsBW3e2JiYQnbdfPsdimkLDgKc5nHJyKyXoO3+t/
S7vpiNxXWOx4hwg9x7fh3So8gKY5+Eq5fw3vbjkXkrsaEkrgO1a1DFifsYB+VQKl
5P6bjAtQvS4nycK/8Xwcqyv4sYUllWKlJtDlLLImxC6NZ+d+5YY77CbT9NnZHYK9
dEyqblqYPimE5VKVoH9/oJdo2MVvJbXpjPOD/LBMxC9/SSX5S8f03XUHWnHkC+P0
XmLKQHo8eUcP3+5Usy1+y5ZhP9b690AAQqFMkypCZWf72pDnaitmrLvTJQ6qz4+K
2KUJjPeHLx/cYj+TH9BTiAAY5T/iAA6wnp+fn3W2hB0XXXdvd9xVynE6LkL1JnFm
TwXW4VroDR/jt3t2EbxFLIz8+6o2xo1kTUezGsMqJcyAP9pRojVxnqQ0FRHJjH/b
KRSE/v94Y+a/AOdBDO5ideGiFdbIUfXSWcDbcVLOEy/bG7FAs8tej1BtFvXIPc/H
98ElHbwzqgllzor/Bhhvq9lpyl486WsYhzArVh9Uf2/sBRepNJLsY3lWYJM3TSEM
7ShKxmnKsRxUhXy4a/hEKSbNArBwU0pCGOuri/yv/tzOFHwE/O2jusgQpR1D6hNp
hLub2ixpe5fSYNspLUseB/e7+wWOoarhCTKBeVU2faqXJ7cUoq9HpaHwzsvS8niN
YCnjKMmROTD5yvnSWLug0taJJfCYAlAb5716IFSpXWFq0wrjplTmETphcyiEc1Yq
Tc+WtpiVZQzUvtBbNOStWHst79P06Ih1E6hR5pLIfMfWdUXIH7o9yS/rXvKebGlu
83ceXHSWySBhEszx+vO49DSNwRNnXxVERaQeXiqGiqS/V4K9eFqPwZce2CRaSMzD
Uk+dJMyov6Q9xiO20eWNqndg/4WTfBv53TKXAMA2tp+VxuTxGq4UcYemtFL42wIV
r1UtS0DwhFK3ZpHsqSyAEzsqWt/U0eBd+mgNGcuHFCK1L+mwM7E53VDUrjMwKPEt
P75kJZcJ0lH/QiD94/hWnp/JGbgoIJoodcWqMqsH8CWMsnCCkOuW7fClYe1flxYK
67CgfwiFxx96nkfpIwMYSqeghpxmD0OjprlUzC/IoWRKZT+7UiRC7O36bWs1//MO
NFvk/fbppb7WKE3bMCzKir3AGik42IYNvAngB17odmMVlmrFQ2po34r6YeY/pdqi
eHXw1RSmbbV/LunAGXkLCRkVPRuJo+uh9IEa8Akn07IlH6KvPoyqBuTiZB2rXYq+
Dnsp0lCynm5zoZdYnqaiOf2sFnTpWWsrsZCdkAyPm7RFHERlMO/Tj6gh/UoZcCBh
FhFOnv4dUEvtRaWVPcNyk8fSR91qnedviluYw9Jsim9aMCog9D8eL01c191Z8L6P
mQyBwF1fgXmxq33gnRLSFgl5x3qX1JiNYxp3+iRfkCUM3lvQ4TuIFNYPLMDG4vis
A+byonajbvRlAUSI4FmSEnXtAhD//AMA8UZLFVSEdWkOPeLjkbV5GdaONpM5ht54
a9uog4Si7Gm8iuQaRD5gzwpHo9f03jS7DGoeKW6/D+WsGdFk88DvPF/VpRAxrFWO
orGYF+sWcb4UWmQeyeTH2nuHPorsmz0Mi6DJDJAUJLiftjAoGv0h/XoLBjzuZTin
SwXZSANyoBO9eNGzToy7Ni8Sg3T5FwAl991g5uTb8giHmky/j4BYC3dGCP+uA4A+
ZfdrBXiND5yI07HsTxx9UCgJ3lG22q3MdjGi13IkL7LH9081/i4kYGWVgOMzX2Ef
hJ/QrgCuiRUjZ2aKeIKqdd/FCRZEdIsWrIo9HmwFhy4=
`pragma protect end_protected
