// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N5AFXHMpvAXLQct+QUgyqwPwAvFsZ0+GR34qPkEhn8RnpdtsYjDAfhdvLsj2lQHE
sHMLffEuhUmkW6nHFapQEdTH8A7hXO49Uq3/sDXq9Wm1jWHlWhtls3+9ue6yv6PA
GCD+ZdfNFB+ymskk6yR2NdBrUFGV1K5e5brk3K7Bmpg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32016)
bzuHCtx8FnBphIRoG1mCu4LXBVcXqTyZsNqroqGE9j47MBIjaaRo8+BwCvb3X5x2
9Gl6xx48Gc8kEcYcZV5stF+pXt+bzqRU6Ovsor0bsgPmF2+pglG+NSQNkSSHDtYA
AXNQWhVT5jT7EGIM79rNyp0uMe00ZtIZmjIVveUxv9hD2+jLp+JZzOA3hT1bGgki
3RUPt6rODdbVZytI8YeFxDWZGEyoiUFvH9YdGx89ZehUlM87yLRvzrndsiSd+NGE
o8MwqBGOrO2ZMC8xouWsMHGI0r3bIR2jFXEnYFZKvID1lYwZRMLtRbyj3/1cwXqO
L/SFFDlP9/QzwhQpKHAUijgYw8T7GwrpffClhzthvfTOw5K5I8Zs4CKTwB4/1abh
JKGyfYV/XiDMPyrpwxGJZWD2IdITSwo9cdv9nqcRZdp81JwgzfdankGP8Y7M2foA
qT6sGK9UldDwmsUvsIdR+85nZBKTx0sOd6aAv/J7IgWP04pHdyRHdFTawFtXX1qi
0xiqpi2F89t1prATGrMlJYZqyq6ZdEQHKDlDhZkRjcXWPL0+s5do/4+dhD+pSktG
B+LzeEJcwVBCe2iVSZVHalLt1TExxGIkrwYNKLdIawn+71MKR/NA/ZWwvagWM+79
+bJUNUIi/px3xnoNhGnvT8N/QgssB/XQUnXKn2IYJb3qGz0xbGvfdYLqhg3boB4A
C/poCFwgQkw3JCozD0RypYT2Zk/Dxs8rS8s8US6TVGuT1jngaWVYT21f+ebSL5zH
arMMAiC50SGlXiDK/ELjy818kZvQfRBcLUm44J1iURu1c3AINWkqNOyYWIkRRDe3
gBVxB5m4doQS0CPUZQM4gJ+VH0p/8FxKgVNx0bS3m9Z6Z+otZxeAmqXfk4v1IHAX
AIMyqNxSzLGNorTk63qV7EI2sZquOLAPJeE0E8Lb4g++MwDZTew1SFwKBSqQTzVg
lKVgTgtm0uVs4fPr+FaliTaCKkGhPNX8qE1T60IOtoz0IBvzE20i2aYUYFk86jOm
SYXhhT1AyhPUC2ALLVDr7WiShPUUnn5kStNFHGXJbjVQ7TmZLqUA4rWMuHcKPMli
gKQ8oqa7vZ5LU9ZDitF3u9Bu5zDnnUHmVZNz+pkj/KlrZ7KVu9cYsH4/soG+1vVC
UhlcRNfYf8kxBJ4icJtwK0i7qOYXA9jNuj1ngXwFBw62fCiCT+TtZyt0hM8HIpxB
gOz8/4HuJql477ja3EoXTQeO1YZeiRdlBF4OSU/u6XU5jxIsJlwsTDX1lqVm+v7w
a3cWxkjq2m4Vg0sJHUEQHSl6DZjgh08SlT4By/IakmwiFSLL5HTZSk72gYRYG7nc
laGRmZns+FRApvgM8H3b3OfBQTn+xbuinf+mm/oo8Scc/YKxA0mPW1X3gEXkNiel
DN37J6svtsvE5eRm9O/T/nC+uGCnrOYCiCYYD1skf/UhqlKzcC68CTBpVXe4Q0Rg
OAZNJYbFjPn5rlx47OhlHEHZgt/PsOVpzTzckqn0DRTHI+YnyCGuJzGfcaNhqA4M
Y5LDYlOWHnCnnBzCeGgZ5WBdgQvgIKgkdc66yUSLpXiuJ3fGh/86JD9PLSy4pM6t
q7k/yQEJZzmuVNeTGWxEvLLWtAP7RIDTHzSS/MZGeKSL7OXde4j3rWd5sN0hNEVR
F8vZN6HOSgPhkrq4d43xhvhgHJYgQF1JNalHQxmB2YuBHZZudZtX09PPLEFcfgQI
XaMb5MUMJIlvaKbULWg8vSG16PWAk3dQj4rcx4uumIXqwbJ0NwdDGGrlKSN/HyHL
eNHp0XfcjK4ldyrRhWNImA5L4/Gh879Uh3vwrfW9S97KP0BAh7Z/P2B5LQO11e4i
8ke3Ox8EA4Snt+8YCyby7wW30k15KQvMqKGRgqhRuGF4j8/8R0S41UeF/7sYOrvP
nZFQS3YjOUG6vDxzsbZDyPiTKJQ0CYCKiHjsWlL5yNE53z+BLP60cqR7dKLSD7ol
ow73nyuHQgEEBMm3H9+Rkyry6k5OX7F5UuNT2VD2NAUFijDMgS/VIV5N5OEBvdY2
kLC1iITj5905FNJet0oE9q1LkaEDuKV7ndf8kw7chxlbjJX9lBbvg1cK0gFoBZWL
t0GURjcXPjVQTZmC5Sx01RQXqs0lqLNUKkV5WR+O+pGZDq5DIhPa5zlKmV1pbKzM
5gHFSTIzq4U+q59+q5H9LUD29KqjCXxw3oR54tDbJLgAQL9Ii0iiWXbbeyej0BWv
M2b3pLmfEgXqhf7/vyzv2t5DAFFzuwLotcFXTJi/JS2BMXyM2qkBncpsnwLg3nge
+QYgokQc4Py7AfkKgmMn07IdVLJngbUQN0VdRNjtSem/HPN8MiNmTCbLf+RqsgMx
yfvi7MDyI+XrLbG2+MeKmSy5T10Slru/MDR9WfDhEym/of9sMsY34uXmCDzInlde
YaoiMXIK12IxBALbBTzZ0rLMhk7Kk4FH7utE+NpHa7kn3Lt8an4NdKeiEcxYQMst
I7Y/D8QqIylqmV5k3gdx5D5/Vx4Y1tnbllzF/2HZdYTvOdA2zLKfp3Ygq7I37cZj
YHgUN2kkksdbYjIvETBdh6u9G4S8kDLPpT39yqNrcJXO1d6wOtpn4udeNG3m+JVp
CzqJnjjQocEi3/bbZ/emS5dFhjsS5OG9RS7BupXkU5qPpBysrMo6dhNt65gB313z
4NS49RySWlzTzamfVZiDkePgIgnEx6uJiUrUvnH3CJ2Ka/8ivb6//+aVJVf95LMG
NP6xJjVya4nVSJ/7pNjjVjMYka1DwolZ1iYtKG7YdnKrUxCzQf8rfvrJCoRH2H7n
LitqR4stniHA6ZAvxyO8DMXRNieEC+zIiq/e3gUjepXZI7hHj2LxP6PEKNsaK9eq
8oExsXrZh64WvEiWbQd7gsUcJ69CFHlx6nKBiONfuuQFPmidY6+O+UZciz0rCPUF
jRxzCQXvU/VCtDK8Lzqiy2KNLEMwtjTBXQO3SsZQXhXZl3J5RJ9/FV6jRIiE7U7V
tWG7QZ/dY2AN70dWMF3CNxezEzRrSq4513S3d1eSQzvaRQIbgjPAp4KrgUKHoUHT
kmpgkOfPkGCkfC2JTBzdpxBVDtVps1O6QbtPnx3TjpGtB9UyJUrYTwqfyAnmwIen
ZBy6NT2NYkAErSTuErOBsrHKBFnp1vCOZ4gjYGiO5mu5Wlx+CHDrX9MyBXJ/AELL
agAHXGnqKbrEfL4YsSTkNuG+iTCVco8vJjRVHogsDYuwHLP3rCjTlBZnEddpUYf/
ldW/T5wrPz+Cdaf3X9kk7TI2npFSeWzZSLoXgT7Py7k/ru256H+AmLfhDYuCj5FG
E0oh7RHX1rQmSRDuRPEt5eir6GPgfGgNvSLBzFEtYK9mmDYS2mMTGLaypZGE6oyO
ffMmIed0CrJr5sLrseVthDlQauRzH6v0WZZWWCU63wyiiPDHX+UH6hRc5OqjRwTG
AHIab4PlesZlbZ+EuKg89tKM9bz/BjCuIBsP/ZVqLdKCl8z9ECRa9Pfe7tVlKlZR
D5kCzT62RdrYUdSHiTdQG7EmrFafwEqUYl1hAVU+G8tgzZ02KviXmcM0FAiWyZ9T
+WgXx5TctCgcBOcqOQ8k+eUur94IFSSue47ULtdOKLVDsR5/uTwRRJ4z5821FVHM
Y+uvWkxM/lNrt6E172UDLx5RSg8SVTqaXuf9ADQYBG5lbTapinXESR6Yt7La98f6
kbw/cKotzFNKdfIjLlS9B0hLlkP5QSgx8ZduH4Ff8zg6LqiPIKEv9tS4hNgxcHrv
6s4VWeet1K/47i+yHpHTTAgQwpeYAgdVx4k/6kcty8c47Pntd5fn383l4WU9BeuS
vEEs4rugom8hdCSD4JGyrKUSwgYBr6p1FmM43DvzXzaqJs+RUty/+uVZaPTgXVHD
kgoxllV4xVA2LXl05wlhB8roO4x6U+7+M65ltJEHUwXww5AjCg3SHCx+slvbMjrC
yuuHq7BTYIbMghvTBpiAoQa0GexgBqMiq5ijboSUCoBPezn45NCFygozKMSJODVq
Yw0xTMzhE+UI1ys1kl/BfJn3+GC5//KqkCZXUibHos3K3KGXf4UlAFNmKgj70Dea
jgsEMVB7smhF+VTIhZqZGXIB8apWgvwu3k5uBiKQ5j0EXq6cLluKchdayG297F73
hlCykTW1Ml1RDJE8hThjf9HdlNUFUhYGQTko8LQG/7+9m2rTzzceKAgub5pr4Eu/
jK5ZElwIY0h/WDaQ7Y9ZIkVXrUl8qdtFY+4ZRIL0HMEdx3nevTvLJVqQ0RPmY6+C
0D9q5n/G9EaRi/Vqo0cLFfyHUc41pxoEBbyLN4LRdN9JlAMt4YJ1I1Wa9XS0eT/p
XD83W6CPNfXep62BEzFS7PUbmgmizYLTIcBdLjdGmkbYLsMxLxy82SaI9Q9wn6Cu
6xwOjqo8XVMbEergxAUTzWMa6whZ66c7SeLt6IQEv7UYRjdhU41lD9BgW0kA3rB5
vR3C5GmtD5MIZ8n7GV/Se+svIv4e9zUBJMZ3Y51jnNLFrKOzIriErK0KMUGvfG/P
Z6ossb69DN9EwmZmQyPMScJLxsh4MaTg4MNlAP+GSjzgytlE5HA30F7VYVRtCDx1
bYBZSxlTUwTjR4dGmCqCKZWNPKz4suXMtnvMHkSGIDErv8TGljpDpXLeeqt3KmN2
8Mht90cVCzjUzdXN7FljoQeTsygfdQZERlhxWT3/ZIbcxdA77597TYlsyGI9xBEq
mXjHm7dtsHc+mF+dsU3d3A75pw1nApjS8r3ZtdLeIT5TUrLthRcMWefC2nnLa//T
5LuSoT2kodKtWVEyxw9KepAKTxGJ+FCGNgi7YYnvbcD2TxdutURuBP+Rak5QxUXz
2Oq/z3/PZ0hLPn2buL2vXeirA2CqQQq2zJp8hPvFhJYa7UCCetIL1c0pGnZxPwRW
8L6/cGImJMPAlrYUsJ8ppURwA5vleQ2Quc755zXGdiMdgx2fUaTxFVpf9nsYd/Zx
fHDQDXHzK2/ElDBqp/DkKRhcKoj14I9S+FyVQ5wCt8evcS730/pAWXmYBjW/72ZN
1hpTzd2nlM+DtCeOAbpMLJ3Zd0XVt2EmBkEDLAWkNyOBlE0kkVT+K4ldpBY8nrUk
i4gV2e99tJExAIs83qq1aOtu13fxIG/CQLH0u4nYnfiurpIOXDWL3I4vVNBOwpLs
qD2mPGJk1JF4pMNKq2Efy6bGljgLznDErPd2dg5ihrn+sd8HFhkgWe64Vqof5Ibx
Weggy1KJcVw79XSQBF2ExuUafok1ZSNM7EdBAVZaYCr4iiwHqjYmfkkjDG12xe0X
CmE9bmuT03PkURdMofzrVf//R/RVtPDULAzaxmHnGm2M3dejNuqM4ax3fU5d1eKm
uCJRGgmg1aXKa5KllZfUIt6gZKtshGMJDPCeBETvzGrAjdGNvKB3nmO09VCxIBCv
OY1jGLxLha5cD5hcZTNg5muLhcvvZ5AHrc3euPefEV3SaGTbJpQCwgprHe0gYapV
0yOcE46zIh7mo3nw3uDAlKhXeJBV7AyBpodXpwdXiWJb02ctjJ4hUxkL1yEdUrQX
Wep1AEpOkcPPQNkVlemP5K4r81IN99pleYaH6aNiiPdMb7hEs0KdB1P3ZGfXMdbL
E2XH4SmXgATE6O+qBoEPF/XM2Q//voLGJcEbOJNkjXkewV3AoQkohDAYPthwszOa
RcnXNE7GEjYe9c8UF9Mqa7PjNWZ0ZU/ucN7p5uTZ5m/urT85YvUDdo9trcBJIqKE
a5HJctjUrTFCvd/9DSdq4rUnQTWsClWijPVzUe0s4Aa0fTbN9VrytuJ3oPQeJQZW
0CZ4hUh59ZbdDkKRPmk6s7DY7aiB+bJx1OvoA605ulCMoIwMsH1F7mAmslAYecov
Q1goa9bXJA1ZWa5nZp3iUanrX3go2z5yTJRc9OV8au370NqpBjcVaIecml4aQDvq
GspA3x3P08QpoqTpBf3HiZo60eq65iQ1QsQ/5dtKuqVYD84s0D9vMzM5JL6kgYeC
JJMoEz/KwGo3OOm9WsTk4QFpRzxjZ/ASX4OHLxLyGltySY7uo3/vb0y/XzHNLCR0
m0D49cJ4wqdzUcPDD+gQ19LrwkDMVGwmOSt7MvsW1MYtA7owpmT+RTXJXebEB6eK
5zTXkOrTJwZBJGfpvW+Sgi/2DAUJ0PF6Wi7l6IU4F8hzBAS7oYLOC31dh40JPvXB
fuvd5j07Y6mPp0XcDHRUCqRvOhMOY15+0T+uXxs0BGtaZfTA/uKY7QdmPjQN0EAS
nQraodNjSTVGMIVvtsu4zej0WgWuRqgIRlqfekYTkkKBdR1euo8O8QGOCrnsRiY5
7k6sytpZurl80VDtBkYowW1ckB4hTG9PUwKrIJxu2zgRSU45962GvirAEZFD1qq6
zQzgDn68fX/7xPZeovcs3yLjXAcOpjPbgvX1pD28pHRaDphNNNNjfnZ4xes+J+bX
k+65P+uTSkQV1o6FPQACsnk81JXh1vL7JjJOvTbnedobE4du4D+H6Qrr9XKyZC/J
euq4szc3lH0nJCW17AVf2l/hrwZzAZEDwelwMsvIE1Z1ctySXTftk58VQ0I4DdLb
CC7Fnsx3ABlnaWhyTpnFOnfOmilgkuOLtqa6VWLd5zb9qcTJ9Wc4LPuLb8lj7MT2
I5i9KSDYPCvwUHWNqUmhwpZTpzgM5/3zI+Fho0NLLVdnqWqPo4hHfIStrl/dMLI6
n20ByJZeKme8uiXYCS3ASXtBz0lv/n3hS+5yL3BuQrr/A1C4fyCJBRgjuC4GRlya
5U7rzo+RIqNA5XlUH5iKIPsASia9YUeKRcBzMZ9lZvhkSmfim7rqZzF81AY8ocq/
SvCoUNUHbY5eySLK+MznJmwGglGrN8mTrFDqAGJ9H2h9acEu9CETxoPFPcuwM+Rd
XMF3Nweexn8qGf5O9rRHv4w6QUjxeMmnx393lwdbDA0MhyExE3RyM8wa/FGBqpd4
t+J0yd7eekLqZ1brdEDsbmZ8yovu+IPTHaKjUCelnmj1YMJMhgK3HRMetiXReLpR
U1KwjUACRYIfpCvIIy0gA40F5R7YdDpEFpkP2N+fqgqjA0SCYU0uVcH4PGs7p10v
8MTuhyFFEpk3ydtyIzzaTiTZ884QXKvimpi5G1XXoDoaeqLj7tfx8lk08Jg694s7
EUi0v2KFIY/lAZsjkGUakEi8QFOkhV6I4fJvxvESasXM8ScpY1WB2IFia0vLY/Dh
QdhiwVGCpWUkDWkl99ZK/abCFpTxeAepvsXdSYR5r0LZzv5T6s0DczNGZwjUB2lp
FUJ93ITwBEFoBMo5My2+e9GrT4ooFghD7Acn7HY9r2ewrtH8tbmWUHoS7nJjTHYc
qGjB3JeGfLMuraapP4sg5rx4CgXF6Of/301twyaA+8FnS9VFRk9Qz3O/kGTjU2jA
+RCB7bCjMVMs/qHFeeFJV1Tb6cFll1DKvvFZ0X4O5TlBNNsIA39EK4dn8EX+OTRZ
mZxRo06v2ouP0j21+pZ+h1HsIWi6N92XbZLZUFL80UNTzDIyMVimoRC6hF4abQqr
yjhanP5YI6thlAc/izkpHkx4r8UeTL+a+LxpHBRky/K6dts/iR9BkCqe/GiZT1B9
Ey1h9zcQ7gleeEMJlm2V1DQDDnr4jqghmdHZmbr7dXKPPNtVSIXYZ6bNwTX9oFeb
LJNacnHUDpcI3kIaKptZdq/Oc5m+10gpWfj+hWh8fsSTeGHGQKuqph5mjkZ6E14x
j97tcFU9Y0K/B/r6cOfTnXJHFkcrbkqBC95GZ8xbTjVTWotPCEXFzeg66vKkeHnw
6YvX+7QfcfHgU3MVH1PDbp1EAgNHIE26wWMpq9jfXM/pX4uUvDkfgwvmOSInx6N8
JMbcPS50LVyp2zw6SJt69OXqoX9+dAQr1qHcaB6U1FJhMTCwB/6HAlkhmMbBjqTZ
nSJJEAzQ9Wlk2SFpH5GZvw3LF3w0/nljEh9P3+IMvMF/rmaMWgUA8d2ENUNbn1Gz
zPji2m7ZsUAqBEofuoke/r1NLx3UCz1/L+XTeBnBt5MVJKxpUovpETfJSdSkG6YU
CUthso3myP2IUlGMr1ExhYGhwCAY59Af3e6DZcoyiTsg6cFhnDqxqlNt5qpjHnaT
RuZbFJUAxgFmf69Azl4DNYLPvy1muZ5UrXjOt9sMu1vWpCUrhfAyaFVDhppUaHia
xm/cCErDbO3EzCA4ClpZBPBnyEhaZRLHjOc+Y7AjFlrTc5MPMuYwzGhZvoMajVys
TjcGLOlyWaPSIJHhTUUkKRSA0fN8G6Lr+pgIPGbKhekQMyeOPZCGj2PBM0HXh28o
DL1lmVxw2uPWXKSIYoDVcpjuRbmH7uZeS3n+IDJAilCGN1J9ghMcHBrwefY+4p5c
rWMAJO2FBmSD7kqB893KTUelLyO6OuA/dSpcMeoYq4de+GYax4jYNKeivFuxsD+q
bQU/d+jRfkGS/ec9Rb2FoNQVTSJBZ3XRyLHt1aeSqZaynaw/zX//g91CP1eTppKa
CG23oEzC75x6EeIGPhucX/rE0JN1OaMWj8LtdZWLku4IejALqw37Xt+T0timBJJ3
xEZO61BaFYq+RiFxaQH5Xs4HNUycYWPevLAFlnvlXvwDgpwjAYFTa+CQGkvsG1vd
iJqeOlXJRVGatJeu1/7K5u/gHNHFyicgieTcYWA08PyM4aeeqVQwB8ovm7wFz5bl
peabISpLK8TtdBlPIfDvZ0NvJcBzwASYbT9jYByax+N251KnkZP4gi6wZMKKPjmc
iDa6y9XwP3KEnGfaAB/1eaXOlkzEJCBW4Hfz0I5x3mDVlEZ0Vb1fkAv31KdPTIIM
hHUhoNkVRIjQs8rbKQGEsR0z8L7Y9meO7OWVbyvt9Fm0DlpFJ8gFGtvVNCwzPd6G
i/ELlA/3/Db9a5B6SLP0XKbFj9pOynFCbvtNxF+6RSMC4AneRbRz1pa6ynivnISD
WKHJRIBxNIRFzMeC9NtKr28yDvaj4SCSD3XO+ZfBbAj9CnrU301oeDapO9EfRKdD
tvwe4n3fEQ6nMGY2s/1EDJGZArBBqS/6b34gqIzeiz8UNJHKc9rbB4Y3EGayDAfV
XKxEcKDax5tMXwdl+b+cyooo5nyP8aCZxvtxEwMLFrUw10s64NRK+fH6q0NJihgq
z1xv1mgicKXH9js5dzjNzo/WDbwA2zGNbyWL+uMCDEs4Qa6QAdvex4fsh+tlJu4i
xLRxxESZHoKFD0zs2lCA5tsXXFQZQ5zUtAeUU+GcCZKuIi3EMLKsGTv6aDRFqZzT
65TzTQwswZrLNWGUfeZBuSy8N9awGM/WL//vx+3xgxYTbtguoV6tVwdNhuJFjlTP
lLdnCm0sPmWn8AgvHVb2M9lqXicmaJpwUFrA6h19TqrK7Ag/fTv6pMtgjsyhESzW
ekntnPU4Wz0KvwC4NVBv6DOBqwzdJn9GQ8iSDmCDEEb1D6GrV4p+EugoGaOxulWH
CxsIoPL01/D9tEgA6OdkMLAyLZq8Nkp3frauk9u7uMHlT0RfRiG/oznZdgF4lxLT
oq0ibotm4hS81F5OFW5x1+Pdway4EzE9MHeM0TMNrSFd5VJHuzPyr5gvEZWeeuo6
RCVIROprpqdpN935l6TDdeXc1SK8UTsCOO4FJtyEyaS02/wrDdYS+TYXGXnrppS5
LbvW4VBPEGCCye7L+KsXhlCPTvZBjilhVq2Ezdnnc+k2BRbiPiNKfBnmlDGQFW/W
hC+zfSwvYcxYWwa5O1NURH7+RBu2j1L+r559nMDdPMaMwgM1AGKixxGLyWXN3Mov
WF9VQvu5GpAMIVoS5EVSpVvQi09ocIgJlcVWGPbkQRkcG21xC/WH/EC98FgyQ4iO
YJPrsqNAYXBLRcFOsF7YYj7Rv8cxWqd9J2fZkSDgOh+t7TUJ7nShbSb4ziuTUnEW
xx8bhm7hoQa45PQyrgeeGH6e6dIj/eZKr7yLlA2Ltzz4p4WGipeN1Hjigpc7g9NM
bNlqkCsgtcpwG7vnaAHAkU8sla7w3jKPi+4GNmvEV9J71f9kGHFMEltTI28w3Asa
tVxbzLqK9zFaqVD9JH5R0brNyDwQShCwpL8hEQITNPLcGGGxyKePcSnGp9AE4SWB
gochOILTOAvgB4ZIkq/7Zov6lZ3KMK86WCBcROkgKClMPq0LkWW8wejmysP6j+Mj
BS4uIV7sBLv2xLsdnyb0i6wQQhyMe9J1unhAOWbKgh6lRncG7bm6RtuuJkMxhcB9
cLR2Vr7MWVdk3xwzo+f+vzbbJYOyro/tX03ewje3g2YP6aFrnTenx/JrfvIZgvvA
aI0gaptce/HSZ1Dif13ngR9ANMavimsJ5P+u07NREny5g3tsBKgTbGbRbJt8hrcg
cbn6MrR0tHWZ4lEZsBUZwKEr0ZCd7BUEzSpVBIsmer3OzktDRzDAxHOtJL/UH3m8
HueQQUHrZGuY+tyLOASQ0Ljx6+U6+VB4o68fMy4phvlYWZCvHDdaq32Xe7KQZJKk
VQ6otR2JqAUtJFY7JYQ50N5uI2iVqkeFypGO6sEWeQtqapOOP2MUdJJjCDTHhN4F
h29rVvgQJ/paTMUJW6kZATeUU+9eBcCM4cue5fMkt23jXUrPR0PVALWfLWzOsjek
1rhNka4ZOpzrd8/5Ax55YCN/mSTtp1LX0GBf/ECO5N9uLEFGpnKxjW48p3UTEijG
uS57DJku+Tzzg+WkzQGWVHA5PTPjNjjlwh4Uaw2hpBFAaQakbuHC9zsVGYDZuP/K
3fVPNb/tttyj+cjRLoQnqt5R/rpCMaWkgI1B+x042ZPhhdRtFsAEd0Ike7tlncvp
FP5SLEMrb8GtIfReIi7RzvtcgK/X8L+2WWvPTPjJaL+IHrMk6TuYph1ZSRO2xMLy
ndTJH5YM2EYnHtJEJ5ypRGMXslR0FmjaQ6lsS4VlHR0FDAw98AV8S1c3XyYUjfmW
3+7YvF1JpfGEf4hqQDTA1YiGl3BOLHXd2huunx2RVxh7us2MUJbVla+F3aBSXWDr
q1xxsDdpCP9z7AyDP2em1658IOgM5UsiiPw8KCadFUNjVxxVC55uOlaQY6gpAg4t
W5X2dtKGVByNeoDpr8pIcEuJtwhTOlhksZWQWAmyM2q+HepL4yKYNUI8Ou14aVAY
mVh7Z4YrWsQKolfDq2PEDqDEFtpuwOxYEdVDDoDL63tRAqicb4439Hqu5pZm/gyo
xTmgLCbIcB0l2hsRwYy6h3RABriowwY4xSbUycwE1OpcgSK5I61WCcdB6Le2MIx6
bs2GEQS5ZEHqAgXqRJMRSP48hWlYgqc6h8XE7AwCqULRxEy4u9Ld6JM1hibbE/C2
qFEu64RkztyQUPrV0LMBd6PqKLe5oJgPPvs2yVQNzlKNMr4C4wDVQRZMUabk/X0+
b1iUzsgqALl4dVr4ZQ7c7rTKzHyNFu2ZuirxlRsfWUne61Ao5QiWo4R1uRtUTSqn
EwkHMJpgh1UGlJ3bxzyZ0n9t0Ib7/r5kJeRFrbRaTupbxNuei1WgME27j4gPqwbX
ApH6Y8wpY1y2apFjT7vyh70PEm6B7qp21BE3ZNZMk0ks8nA6B1TGXj+VW4KibtM5
JrAbbqxoc17yZkwYpB9P8h1zNF35juS0SSo4DRVLZMyRm9zEprHClkEEpcWZPssd
sYfJs6JQmzVIF3dG9Qv2Yp/A6YzduDkdziw31SteVV+2EZL3I5mJToBnqvsi71r0
QpXsyKE/poEC7j2YaquzEBxJOSrHtPteX8guH9TO0VjRHuOthAww9dXUxLiD4JEU
hmT4e1JqgQSyVqC7Dom3Uue20J1YCqyr4Pj4jS4qBBimOOuQwTyvsgrdBFS0cLNH
F0m2488pLPJNozltth//81Ubs2hXJbDumQmG7FVt5SMpWqvqPQ5UIYXpExVsL+LS
AHF/BczPGGq5o6n6dDptcOcFkEAh8rIUdjF9pGjPpvD8cGot3KRtrNO3DDnHghh3
WCa7eHXSCcJTcpEdKruxUzsKMsh1D2KzFANAxgemRTJX9mWigGorASV9EvFEXEkJ
tQlnXsh+37rtWIeec0aOuwSW8FzCYWXi41KSjSodfQe2OiQhfK2Qpv5itU5CvLlW
x4RyctlY35tMNT4iahKApzldkf+uAoPRLJ+jNSNYC98e11qASgs8KLaj56U8fipm
6O9ALq+H7VP+Asa2D1pUdl1Dl/AocGme4VqL9RkI98MhEgaVN+kPwC9l1CG+yxE8
/VfoGUxL9lK04iQxdnjgL/bql07v8VCpW6i9k0arhysdWkVy2ranZM0qT32pAQ7i
RIjYzId+ZXQtgjGwc/Q8hTnsPC4mmt861W3JJFqAikzze11WnMFPEy4dkbcOcEQ6
QTEFDF8sxJXeaNIKNvc8mEu9zHTbYlvgaw1JX/4H7B/Pl+UHHbKxd/NeOiEKexmj
APhPR8WLyq4JxIrNXamH7zITDInSzVV9ggtHaShOAvqD+JmFT4/fsCj3pC5FM2xy
w6i0m9W//9U0mg9d80eDN5yIqw/0D8Ths6repxbOydxF4IgbREmJWMmQNQCV8JCs
EP2etjEk3jXR5yRzCmLbV6fuznDrtHP3qPPJWGMza9RNf5IsuTf7IY4Ezocca6Bn
hhOwbORnn2/ghW6ZjAXbCeZNRd/h3gnigdkGl/Z4YlB3+8z7l9jpZPu6/m0HnMD4
Wknc9dkNotGTIqbW7/EbZ8lF7Z4foC3YxwB4foMASCiNkfdMAHpxdayH/1cYeTVq
WjpP51rYPdUBBSFhr083HWQ4PWMTdv2fLiVJiIkMko33dx/dG5uTO3rLCUtoY3DP
jOEuovt4p9fkugCva38RS77j0LpAjRUGmpWpi9ZcTzSWHes8S+J/WDzup2T6duh5
tz2MMXNbVuh71Cooqgvg1wfRwIR3BXNg2F8+vkpGh1gwautvffc07/oC+TWHbfqa
t1+aZEO2juLZnZsx1TpTor2eXHrbv7SIc6SVsDmF7QnWqN3Qe7fpX/y7BLFxOA9j
FgpaiijE8f7zTeCY2W44MCsNj95WWIg4xvSLas1Ja3rCZOTQzSFhcKk6NntDoD7V
0ujFl3VRrJeZ+v9IiNOA+HNA+ynsu8LY1pTN4h2KOtJePNv5nESCiZ12XfDeUbzi
Y2gIke6gAVj/JoTYGnodLXPVySit1CbuFSJu8nJrEWUqSKTkFHr9xAnuGOYJj1fd
woM8GS0vQMncB9vLi07JMoe+Rm5H4yvagfWK5XOsqqurotRYm+QKHtLgmDlVNiXy
RRtio20AjGCCRD3A/EWVZh3Pd/3oNy2V8Bq5CASyyjh8u7rbQ243bhJOGL8iXzTN
zKotFtNHYchzmkEundjUjCqXrlGJ52VlCIlHXINxcNoTv/fnQeL1Tvw6y5Prz0NG
M0xWCLiAKgAKLpPw7DirBTGFICZKDVR7VA76cRnKIa0MG2KQrGH+OMY2NOiMoJ94
4xY6cum2oUUBW7FsnfkclK8OQgRDEUz6wvegd1N21rh+IZjobjSxrlODYZBfZUGz
dnGbREntnkBp2hcI2DTcrcBIbeJN5iYEwJFjm+Fp5TB8rapr294L8Vna7BklsCU0
E7801UOZA6ywH+nKivJkBJerxi0VuQQOMI24UFpZg7mhyxpP/HRZ5pu1BBWQSswK
2r1YWIi1g6hRxmxiJgrW5TSw5BBQVdeiabR9BGzakjTuriMZixChS5vGns2akL7g
cvbn5D0ZmUC0SVL4X4avKbZwpRVRvsXENZSFuKq/hIJBhdV8VEfXu8Plq6FaoCeo
qeMhVjZ4EUYBXLuh71IDx2reyn76u84IkcPtE4BKZW/PbMYBtWDLxHz8bnphBA4k
3aoBf/i9wvY/1Aeiwt29UTy6CDnepITBjE4yh51sqTcETaMdGLhz38i8lwU0BWQf
q0qbcLQB+zS2t2YmXJq4cLVzT8VSczhjKUjqZN55efmpLMuc8lssOjFUzg3WiRf1
HY5wmsGmgVcx0ldo88zu2efm05Kz1Ik4P8EYxMsecqHnpQbaPrWSpQRtl5tNDCQJ
N/3Fx6axH1Tfz+GBtYtImtWuNI+poABtZnHgkpnuuArw1VjEPVEZKmr3dB86NMYq
rXtoA8cWX/fIcLW+ud1e9mN2ZmCO2Pq3CfOtl5fJHweSesapgezkUBsm8QsAklPN
yNv+xzvunyJonFgEdJUQZgZoMzmmxjDrIMIuuG0NofxcCbCa3Fi0ZmYc0CWUAKbv
avPz7vRVdKrQNK7wXR8mRhT7MZqZQ7Svz1DPVT+WzMjIsVM+/BjZAGT9DDJ/F/pJ
g83UjILapNEXUFC94sVqWvVSaqObqt5shIVUd2WQF4r5jBNWtIgfzzei7c/PCK6l
q4pWH5p50bFJYtif+QWVCLF4CS9pwdCm2R8G6U8WNEu0sNdBpf4TnsgiftIvxCXc
sWYKzztLj6vho4FhmQCfkypZ5SUjkTXd7F1WpHXlLEehPuPy+eEhVGY9nM+lYUk4
aaeBhVB1AVoVG6kdsKBGya+x4iM5NacRaoJbBat2IltaoDm2d8ngKpS2bjLjNh7d
p0OZQ3hQmcR8NzaKHM4HBD5EFVbjOSmoq6HDf3CqAHu5PN2VOus0VvUPE8zJRMQr
gDnYMovbpRLUmTeUvHTHrNcwDd0Ij39aWtTKdOAZugCYxmOvD+fR0QzHhqH83l5a
s6MkJLVWRUO9PWrG+VEtynYQaYAWSB1599oYUQAm8MoP9WtwQMOkXJSLkw+pgTCB
TeYbcB5PyNYf2cW9fqaH6SunNXAD0zGmyZna0l+TlL09NuQIBUCYPAY2jzp5in1+
BdplPIHSjSWMS33aPYky/TKGC517y4NBIh+x1KlXVZAuH+tLB1OOEW73IEdhsopo
6ro628euG3/a5kAJjuQS8MoByj5uV5mUePacT5+JmCsdD62IMz2R62mF1AITvdhw
e+IMpfl+4pjfd2eOVWyVkKBhAraFcLFv6zo1Nv4ippHOQ9hir1W7qbU2dmwTndTn
VQccvhHvHdWIQpchXIVONgTTuilRVFrXwsojQsDYQLkNF6U0EOz0lvEdjaZ4mlku
fprrILOWWL84BfGNWSuAZ8lcpKDNrxFdfAKDl0TjTF8JWUBI6qAsfkFvkkSGhLed
fCyOwCavhOYb/0OTJGjUsdDPm2Gk79BxG12jVDRGT5YKVDHfrGdfRx3hTj+T2Rdi
/0BOLEovlPj3cY3jGARe0+Y74NHPknBt8/udfwnj09x1loOMeP9rIJh3vM6vyUMG
Lqz+teJyWTVBeb222VoaMw6aX15eNNmroPRh5+Hl/NZkbGSSiqRwGpTUsd9l5j6g
vuZdCA4lmj+eFaR+PJycBmZuoFtGhx6A4PP2nP/nIQsyV6JxnH+eOwCpf+oD060V
2fqn1svhfdL6XDA54VXtS1qtn576UZjg80j+wis7yDaRivvtUYNEf4W41X93mUUU
4KsMk63ktzB5LeYSa1dhGxbHdndqIQ2rTWnNx10ruBq6Dp3+yrwi35QSGIi78mXg
a9b4QeKr3OzR9BbTKR6mUE+1IHTTJeGNW/Fj16Z7kXfgoxIA7kSiAPP6xqQ9ZUQe
k3xwGW5/WwuWov91NyXnks5Sfun/O0k9RJpSBivvZkZYVxCwlVLUeZlf21ID46mS
lmvXL8BQAUvPrtSRBmo8E4tYcjOfb4lmO0KdUqjvW8WwNwaA5XfpUpLSyN80KYvi
xtm7A0DK/B3xdVc+z6bOmxbrzatw77IwaV5KIhWS0sjT76MkTZWwORXgxhW7MyKg
hg2VYJkLfJGLXn/angdt674te8dEhZ8X5z8d2eLErsU7+pOPYBasPc3+BStSTGIf
38V8hPhHx1LRakIfyTFjY9w0qzwn/BKCm+/oSznS8pLJ3xO65/EXFTwtxRR433/T
SazQ9hO+SKNdxotxRwx3EuRXtRb/ovgxVUqGMlBkJqgnQl0RuR83Rsak4iSUtdBi
LWRiX9yxjdjlVl8iFF4+cCshwydeAQKAYa4/Z/89+dqze7Qk9qdDZ4X7lESbanTL
aTjJC8Jt/ROxLSArQa145iEyXxogi1YOeShXnZ0yqb2IW9bp43PBtZoFDlFRidhJ
H3vWH6Y9xU4EFEhjIT8fcs4haKZUWy6A5x07lz5DRXLo9++nL6kAoXMB/Vl4krLR
2GX+hc8ZEYebib/OlV4Fx8r9LHswLboYvsVLVRMIKCNcIKuH7rwyl1eoTHDZ6SkI
NITV7DlzfuWm03ZvIrG14d7nxjW/k8D0e8sEmy+qV4JXx0HWrl7fqPu1oV1ZyHeL
4OtZuY+IynLqlQFeNjpC9zGsFGYwvQZCSWfftTjR0sNLxEFTemSiMsM9ZCzHzyxr
T4FJf0CrSMsyWVcxRLDqyh/zImlXZ4GW05leQNgCAG8KbQrrn0BYTJT6tfTvzBoT
/+mcFWEM601vGfOoQkMcZfV32vvZtIfe9Urfwq3WCqL/IRALbUPvbFx/YoklIeyD
/ZMT9ljI01lW0DfCTuZsmamOr5kz0X9EK3Pb5O/sv+KO02vreeZj8o1ZWo6oyJST
7YrDRlJ+y0ONig/MxDN8HJeQBBwBIjsO0vHfUBwJpQX9J4ABsG6RbfnRwJwER77F
418DnmT6IlWMoe81XDM+dGAcJXeQCmdH91fxjAGfB/oQejaWELj8/OLBn2gMSDcR
BQCzYbBAfgtNZ8m4jf7gN1cgkb5w2Pf9q+ryV91j1vt4efBRSJA0K6iVOBuVv4+F
a4qlWVTjXkkQN9CI/vRBEQF7N/MJON08AreT2UDogRVBD+bGu8ew5AMFMEmjMkck
TCiiyfEGcFfySFJCiCb7FgctCOejf9R6oANqrNhEuOUDb+EjqkEuLdfyEVRhe/Dw
G2n2KAmD0PPJ+RgFPxwRqDXhKYYGMWhtmktHtWlBob3XwbZ+3jiJhxJZHu75L3G1
9OHh7GzjMwfFDWma2gEvtLTa8zsGLjMgrQqqUSwQ74CJcLeXa006+M39Q+Qk63jU
lzl5o8RVGF9Ob1yIjD/e2OCbSQIoqN3D8ehAEV6A0FiTZaApcC3Gn3FAszchMobO
8rKsM6W4qNGWq8wXkKiy+aj6YQ4QuuAXtU9vGtRUWmA1Uc9GrX96xVJdm/tZRLM2
F/ZLoVN1aHvlDnd2zZ82CpVtHYhlxK/K0oFrshq2Q3iywaMVDA3KWGbX5dA2+Ntn
/k1GRp/sE2gxhDGX2Cyv1hozxZ6N/kU2mrzh69sEaJW+C7aq2kNLFv+4KlmKUTPu
nd9gDVHxY2HMszniR+9FnR76TMP9/xYBeSvikzc8F3ydFoINB69RtN7PJFNZHZYV
EPfnAmKU8OidZIcXEhnede+ay4SYVA6mmGh/slGxoac0euFYSZYAABuNyeNluz8u
TpOfVwgycVdnCL10hyfLzlMYUY55pa9MlRZZS+qOJAsppZ4WnJA5e8SL1ywbJAXl
EprEe33FwluKvHHz/mkSFG3vRfNiysBkz5jpt8jXOhhSfITpulQpGDxOdWbjSXUO
evVHtMTf9j49fHiystOAnA8GVHrpgxtUKHp/e7xbEEdCFejwFtjyb4BWOeDVgnbP
IQnzAhjwj7c/uHZqEcADozya1BFs82rI0orUcYAt1q5i0jVMncFUHZQSpPG2oeko
00gh+mYRmc9sMKHK/W5ArS6N3BNE9T/VFgJYlrlqbYQGRuhjjub2k+/Mjtit0InC
Tx0uiFOCd4iz+YDm0NBX9uols8J/TpQRnDFjjQlLnGtlfvmeLu6mLjVHjjWM/2Y0
XiZBk5k1oSSO0JKPARt4f27OAGe9sP5uEXXWzv6RMgtimLq1y2ZrXUX+OCXDko5b
W4LC0ewBEbC6AozerN01Mah2kCOzex2qhzSjCO8MHHtX2WiDsv8mWEUOnlZ9r1uy
lxuJRfLSA90+LbDppAlOIWeHFTWc0HzH1gvAcpUT1uZLBIfpnfaypyP1OO3t2TRn
A5RqBH+HCysz6xepnla3DnK7lWlpwbp/m+CDrH62Zc+W1ZEb4HC68I5Yygq3HjF3
HY2qlQMu+er3vxZC9gYLP/fkUFQjZePP4qqILD/wYFExq+8JOndHcCSkQM9N7FLS
8m0F+okNYRjIHwhs+SC6IH0MVVDBMFdQZjByEzB50kgGwXSspJqVeVUPt9mnIcKo
YGZ08dE5kNfNVU8MlveblJXWr0gbQD1H9wwB9jzXGHnXjdMV96SP46nLOQTkh9dw
QYiLfUbhxOWrsMyNZiC/fZcwwt17oNf1g9vUQ2XK7m01k39w0nVrK2k9ZY9jRcBZ
8vUS9gcfxxg43mKsamnQvDHxTkzWM6cpBiszBDFmH061b9UC5vGR7LTYudo69RbP
EiZgGZKG1pFGPoAfZTbuZF6LR6Wr7pa0yZ4BBsD6eNmQAtuMFisen1LNQj9xYhTf
83FB0lLdjnKmjjF5f8HwHz3FqFnNCHPVABPUw0nv/6Evz/yCEESMa4jsk1vSZwOw
ZadDxtS/7MPhJndxSfqlgWZGAvGQYEhwfN1/JgN6kGr1SBw00Pgci7YZMfB20tem
TL5ha3rV+xunhNuge8IJhHbwY43xPi+ShCLSufmQru1vKXwitpOyYdmyfdylFJjB
dlY6zbLYOUEkiyGMdbj6qGhC59ywa2ikXit4+TS/q0IzEkXCnokvYO29wcApbTAC
/n6EB2aTUSGVS7FNnU9/zBzOygfz3YQ1RjZB3UTkfqmEsgEMK09yYlyhu8/hs2xh
MsnQGwEk/49JBM/Vxco6zhLG5zpRjhe0vLLEmlL6dh7RJS7D9nSzezlTDG72Nv+N
zzfMWcmucHwu0YWCFfe8MXB4e40m4pRuiXlWPhHrWWW9lSnGF7CmqBXcPhALDAwh
dkZMiJ5ojtfKoK6ZLIoeB22MsLpb62YhK6jz5D0dHALrGf6m8v8t3JU0EllGO2VF
Zq2eZMEj7mvjez40EV/gas8e0OUVzNpeYV4UsJ1hJ41mC7EN3O5MIelDUGfAhJ2c
VL3F4gVfMXBXUNvjAlwnr5hIRoYAMTdXOu+blVrloAEqb+l0GhvP7kSpQtU9OLsD
LD8nbW3XQUgTvr8QPPupylD3Dbs7R9ah71Kovj6158o5Zbke2voDWcy7nfYBNSRj
SRNr3cAnxFuhUaYqbjdm2/WQ3DhD8mBFKshuijBsNmsX+KLgxmgeHdzKQvt5hBF+
eAZqvEXHEzvmAu0Y+b/pSIm/6Bv6Ht/4PzePged5dBwdeziSTvaaWlzwGBhKrbsu
Fg9wcj/JXoP4t+D8WEYQFvFMlrmttU6bsRP9h1nvx/omNT6RkR0W6iM+1yKbHsAL
5n4WKg3cLYfUOoNuS+hmVL+0ONSqUaybCm4x7CCIPenO0dUTxhPhyWEgLgN/oNmX
PAEBnOBR+Fsio07fAClCDLSwLdREjWFe37V/R2dm3rrr0t69LZ4qfl8hKlohPA9O
cumnIhl9o5wC99D/RRUrCNsaVuNzbmP3Gic1pdREB3+kKkzO1Z5hSNQtu8gEIU2D
8SDGXMbetVu9TTNCoJnJLrGWnKaotKeMCYdtsqCw5fHPC1C+bdd8Jg2xVSYICM8q
6lmtMw19prRaZlZSeEUK6xL0svbfvwaA5FjQSVgeDwKt/hGS02Evk2SIMkb73mMC
XpXrMD/uj9Ra87L/jCLe263iOfmCSJeS7KRMnizSvrBQhfkZ67kPIeVI3ncp7bi9
9G3jjUW5I03mqP77/1IQlzsDYqZ657qK5rAo0lU1ukVQy017AMVV1bqevRVSdFyE
JdNydg2a+UlJMt5Jrpu80Gz+Y3wDtWFqf3Q7JDkOAfey8mRd29wAd0s6gLI9Wu1q
nuGl3N/OZyJTE4qeUa8xI0y85o74XujjgOa2Wp1Q3O5XHsgWULJPzYSn/IAm3WE5
1sBQ5SbP4U7FhV6M12ik1RBgudlwY2x/X53EQMceSO7LVHoeMUD7XfwPR6jMCWVh
kgLow+H13xLSS1MbX5bwMcEnZaXXHXGMF9+XrbqTjjMdK9JisB+2rrXMGvCBTUKP
EPBe+pfMAfhQqEUriJB4CUNpccnETralmcekPMv2uCPFlj4PhyYLdC7+j+KTM127
nA6Hlms9jw9m2hinNF8mgQiPVoksk39gWXIyY3nUKkgaLrhsKJm6WqQnqSZykGrt
vGCPC3eUnGi1WzkuFi7tysL9J5mH2cxCpeL4dI8EJVWRmRuebjDS+f5KRw+a94BB
4DwlnFp+UWeszmL6ew0nK6hgPK/+/HUPmq4goz9YvO/u/ciYflEnd9Rd6F13xgOh
ouJqntKFhP/mayanhblSPDMp031EIRm08hJOs67KeE5ROnWN37JxGR5i81ndQrbx
zd1o6k4AENZxKOkdpGT7YsTUSBIfapag8en91E/xfklEThZ+8Qb7Nw4mUnpzek4v
vQHuUuKWDxQ0fypPj65h42mAAT7n7Djtz5HrAcuHzKOPyEEo/p1ungpozI18IV9b
c1eoKroTnKFK7P8oK/tcP2F/0GFZ7ymlp9uG2C6KRXeP7gbbRK/DsN6sqY8uHHZy
Fd/e2BT5nx9ctbsNddUBPRUCYhHxuvjJm6Hivx52S0gzBDD3kdV2wj3mKDTsMoYV
RLI8QSOtcPJ/mpNZ1PQzPUP1xhXW4Yw8s2sys5yiiu1odyjucCp//AVmrLVPxkFc
baR+WAo5g3V2GnKbcqs7SAuRP7DRMtK044I8jucjt8k7EeqkJTNm2emS7pKgAAiN
UdluAqOq1I0NL0Y0kJL3HlQ3lWwIHMV4Y4tFdo1yvKJeZuz3Z4MHNaXhGd88KTr9
ndcw9Nx8Omj8jABTENMKoHT27oMozCbtEUiyCWb0eJUTcVgWGdS+c71pGCNtsmG+
ZVJ62hpdUtPEXvl93Ht5ii2tJVErYovDa3BnR/ICwibeDCdgTdEYj+tJ997rFE4k
F0LN4/rWYKTfpvQiPrOMZEk0EBHxEL34+gmj14xFSM5v3w7hoNQyOwcNzkng7DPq
nT+cDO0wTeGMQH5zCZnr83Y9n2kZlzDNRQqkncNjFkuyo3q9gxl6FaV/WU9+iXSv
tMp5dSWnEKfUoRuwNZCMAAOYc7nYz6epbQn6oHCbcDQY94KtOdDJPOPcccCJviXh
5Fy/urBvncHD6CoywUBRr3eRMHzAJJIU0QiROUfv2lU7AsL4HTQsPnrhkQLP3D5m
YFDWTjAMLh2E0dn6BpzR9alg1QuVK6AV7nIV3QlloZEYoeOErxXTfANmfIBfjs4T
otP8Oj2hW2Bxkp6X//7nZSWSPB3wC0LU+BoYqMSIuloqR8iebBXZ52dTsthzZJiQ
DvGtEhqsTyFXAufDnU/qogjQvz99ThsADCEuV++0InJTJ/kfKhBIRmmycc+66wCk
SKRL5LrHqJUwJbvgqglU1BYGlxxF4rYWgyRGid9IYOgbP7cG/wFwSB6QQ5sndLU5
0JxpCDnBwmn0HbNEjFIPxcb4LgvQht9+eoIT2uU3+Y3E4hpc21FqjcJvplKthv4v
mDyn4xIOTuinf5WOcEKJvU7uWEQgltRw/nrelgOClgikJZ6srQBgUvxv6LL9H5U+
79TvowLt63HFUX0PItNTnGlbNnowgGVX7ph+0rDn2iupkqWutLzYJR0Gr/VHfZRl
zLdNPb6V2TyxWHLA7HyIEdJEveEwuewHqAx8ZVxFK2s8exH9GviJAe4//+Zl0UNd
hsvtsKfQeJY1dcEad8Fe1dbDztp+RnNTO1BG6vFO/cefKxXSixfkSjJkOessqTPj
k5TUBJuZTSki7AUB3QL3KewQQroWoNlyCN4nfMThut4Vk1bZwk2JKbvrMA4PeRtg
EBBpddvkWB2s+o0SB79FqiXrE1yYgmu/vgk2jJphPXsky3PtTQ6RiyRo8US6YeZO
LwkjNuKpgo0MZbwXNKnHADmgdYabQmG543ka/GePDXnVC/icN81supKnDX/eEGvm
dqmrCR/Iz9twqNEEpJHPAaSBSi6Isz/fqSyWKBtbq1X8Zbe+OLWC2oNKKgS8L3N+
6Hwqd77AZ+8fQvhUAdBY8MzbXEIIKrTTwFzwxlr9KQx4pXUmHENainHf8S8Y78lx
UT6uRRq0traawPnKu+9jWoqNRFvorA9V+OWghpxIrxbAsIE1WPdTfv5zKnMEr5qv
Xi5JQgech7noYh09+jS2hdK4SMm/VkfEPP8267T7MJdqQOOe3sPhaj/4/EDd/3Wd
sWZu71H4b2xTYyvr0l1E5sXyQU/3cwwQHasBVFs7pUZoJVieznZNBZbAb6/Pj6w6
VtEpoCMmsXMqsOL5elBM31NbRU/GipYdfEXbzCH5ursiaAVAAavkA0kLidH/cAYd
renrRWnLlTNk6aCAlFOPb462zWks4doGVpYgNgxwe/zGYaXgWoATXy7TKkBKTIfF
Osi3NILOuiyOOvuszPk6G6XHV+Sp8I5MyL8i37AOggEir9210cP46EWQOAkjymB1
Cft5KLUSt55XwJU8JGgjwsEDqM+VDICc/APD5UJcy2iv25ygFn0tPr06o7HULCu5
m8VJtdKh6ecvlva4sWN+mzxlXY6Qs377OUZDI5qfJKpZxWdYQhQU3Xmu87eR19nj
NmOd0hBMWXtn68yphToP3cVGPuhHj/XtutL5wH/P61FieAVsFb5h5bURpiCiNoHn
uEnR+cxmIHhlNd002MLZmtG5vMoNX9yYlYZov922AxFjlE84ZEEOz8Ln4GvQ+DWo
Z8p+UANHZ0dPrmxAEKQnmWjIeIeVLOFuxULkuW71slZ2PjUakj/gU2ldAuE7SSZ2
ezJ1fKkjQUzXTwJNiGeTWz9VcM0pv0n1JF6NjvLFQB22jHEOWF14ZcT2TitFq5Nc
5sKFZjcERdDJuZgX1yY0wFV74XU1L8A5zw2H6OiWzPiMorT7mUpVvvhcVsNdcGkJ
ZrzWuBSrs/dHx4Q0Y8ILvTg1Qt9GR6MCBk4sg9NnoeuYML7dra6Nh1dLe0zzb53y
SbNfX6dsZ/4NO//3BlHtm4VNSIVRH9DnU5hFQIhqLxv1F3IpdPz8/z/Xjr5/mU82
AeoIYRTDZqTI/I3lYY/FPoyejFdG8qaXtzhgNievlVZTLlrEFgo5wguulLshtUeE
22k1KwalInmNPBsaYMhBL4Gshrg1mMhrqitTwyTjNHOoKNraFS3qmFlZ9uxdHQFB
KCq9D6HKHqIwTZ0pOGxBpwEaQyOv4oUbcceRhd7WkRdsy0rOOPjbboelgQAhq/pK
0OrEQ3FAaq6whLV8nTZHZPWeLrjTSg8oZ2ijW+ACux53oVgq9zCnn1MO/1Zsu9sI
3MDp58Xlc90VPW3sPdmch82VWJfqvmusBulHwlmKkdeu7JFkjjTdSLYUjM0JUeZ5
Sl97XBkXQqxLGoezvNzHzIYJ9FHAYIIcyagkdMm/UTT6/rR0uCEYhlYphYepEIXq
GreeB61rikWKn2o624brd0jBIFkWDHTeoMOp5inBhxyIl0YGoIDvTCIL3wKQvGi7
OVuz92OjpOjCR3qCmUjgRPpu2xLAKHMeZJSry4iapS3/P8jR/lAJ3LZ4Fr4UG9LN
oVh/P+OXTtiei/6gNfBwDroJVzPFBGICf9G7NK+e9Hpyyf2BASFvbpCWJ/e4PPoJ
dLnsJKSPizBrXUy9IlBp/acacpsXOFvxvKQHImGxiXq198hW4WJzyiJd39Vq+0j9
x903p6j0jQNzbXwKR8DCcUXtFQKs1488VOmUFNssESDLZhtdmxtS75bXrf02Krbe
JIFUBXz8j38rVnCtigQUlNCYXwk+A32eHB4rlzpc8b53E/wpYVRVXcZ/4HFd1hq/
Is1Hy3N2cosP+CsmGCngHUgcQloRgycZTiiOnFtumsf6IqJx/v/zaYJE2SL3RoHr
by+6kIACfTm4g0+/zE0rZeukSxzR860oFggNrCd4s/+MfS3w6qOW6ufCrdfjiHTP
Cis4ioVOFQ553Pdx0v5QZZduSSayfrjHrtXSxgdse6PXqZhcIi3iWBsthAuh4EgP
Kae4p+/rlZyxM5P/HRX3s+dipoW5pFb0GppcLxIgfXeegzVhtVCt72Ky0Zx5O7lp
NMsjFpku1ZasWvrznAfGC/4zo0om4s64blIAa54Om8ATgdwQqLLMjKrtLpFAc1G1
IGS1FpDsibn3qH3S5vn9+56cYEIzinSJJhekM56hJEygi+FQTeVVtG6KORXedP5y
kNw+dq4dRKL4ZGwiK234k1fUzhc9sBqvVkitTvj2/zhT+Rhwm6DQfUSZXiiCPhsA
toOW6OPXnqkSh3EU2WbOjv3I4VGKXnGjouU6V166f2IiUptINVshnx4ynxPg7cON
arssGpb/LqBT8HxQzqLjhxtYkof1E/fWwBFO9jyLqtb884V/Fw03g/ohcsQ31ga/
uJnMdxb6hSmMshaLmAinCI2Hl9F4gBzO8LZwe4PnG5mofD8uUgEY29Pb8R4aHNvx
odhn9MPlXRssYqqnWhjwCtEBjCpaP71TtBYEpbyumyZcNDUIauV9fJYIyTDsbCoU
MxCw4VTivxDp9HM+Z1zy7ZK7DAITb+O4eJvEbcVPzHLmY3fxMfd8wgE84Tg6z1wj
ukUYOprfpKAifrCIWc/sNo+unpgL4E9vaDNUBGa4sGmnhurIJEDTS/US6iQFmSlW
x6IN60GFdPh1AhrP8zlBNlqukLWvCqDQxwppUluU9EDKprXfHMAu8rFyq7csHhs/
aq2mjlX4MC5h1MTNF4RUO9xyiwIf3wdwBOsGZLQkx92H1DnC84x2NAbEmt91YzzZ
DUq0Z9dG4isul/eN2Gw2SEjiiw00wt+Hz1L4LRARdMKViQMT5U7X58+u/szWbA03
E6VR9NtUyLluS9fwS5FCXK9b6zV7fWpiVVvsnREdVU9VU9E3CXdj3fj6HmOC9p7M
FJvChenIOGWCuRTSLmamFcHBVblg5yu9mna7NLoE6FR/OOR3zTwxYZkQjjQ6Av4B
2vT3Ph2ybdsCCqIUquUIAU8oJTYOKzpN9f2Uy3EeB+gZSIZMU4lNGwk7BiAazBFH
86HMUQ/WaMhMSsNQcp/YbJ/b4m31BTd8lCGwxFbzGvn7p5M1C6w2EspJsTNcGb75
p8KmFpmigtbHweBZbPHXRjsy6hO4onugdN0+/4dTYA1FOh9vK1fgte2R8TXXmBOs
jDwrAZy0jAddXLaNQFH6O+ONwPwfkFE/KwgfjqZkmZ3S5BYwKpRMWmOUaX6urAlr
qJmVx02YpN9G1WJjEt7LXKr+H9qG6WmRq2ZiEjMwEzbQzqaMj3Z3zZ1vxyQwfKD2
vqMdJA65Eqiia/olKjTmVxtSHGl8nTQjRDNBuUZYLsm1qqnaQr5ziz+9L6Tu1J4k
UsiDnYkdifP8TZ8ZlwkqLALlh6/A4avvDui3L4lZ9vomIe/1ooF95Hgm0Yo0d8yb
RBqghyTCo83/GQICZy2NyDEmfdAdAQitS9TICqoNEuplCkWKT1pnLuo0mCQ5XJy/
JmwzzeLoir0QF6ZmBBO6c0wx/01G9TLBAOmkgA1OVI+lkgp7g2tsSmEe63eBB9iI
m8+gUB6nkVT8pNVF6/euqJZHtLXF3SeJEtnKyaWPQUi4Z536cf8YTKfdyVBFbpDt
17CXPwG333vi0vYJKAmdRJljQD3xgXijBTZV473mLkYilYgtECLexKJk2/CwtesJ
hkhWhRYseDVUpnExpgcFOOpcfUAktVicyDIaIQ21r+KmmIIn3swhBx3kO6w15xW+
oIcOPK2AGKEWYIugj7XE6UUPR9a0oWExyK5+USgPuDTu2aCJhrBIAGi3SspqHvSE
5J66i7PmJtnovr5exp49sZYTvFsiDnAvVirDR/Uhb0vC+cuhrUghXs30Nt9iHzwF
9RkS92zShMZl7NuzT9VJyuiS/qLyWRgimbay5eXzHsOBIa7YgkxibjWoOmmMRkta
DrnoFWJIiYU/3xF+NovFofrHS2tiycqxRlFzSVh3xictbID+riRpZV5sI1tpFPOG
u+15W8ani96xnk44sLHLUxTJWhrH0jwuhcjdHqtB2HoTlGfkME1qcsKrM7tgMD37
FRiYOeolOzLGewhgAS9qzoq1008FRIb352bvN8gIJFboTpMwZL6ZGwOkLclri6tZ
P7AgX0xY18Dcsxuf6v+MOtAv5wiYAxzfIwIf5WC7TllJ/v4QP5NPiw3kVKYi75JF
7TLFtilvDwjybnYxxGZP5apB1nTGQaxfqiwAEOED07iUb32BcG8G5CXqVXbQu5yw
5dAtQ361LK1QKRtRuXdu48tU/ROOD2t20Tgc4CjtB+wkyOEHPP34+sv8+cLcGgK6
y0hyDTXphH0mwTWinUd7enCECivA6+YWiI2jwFH4UhiMQVOSF67qyyYZgK+S3+Ga
v+8Bt9SZk/myxmWh30sRu6pbNq5Jc8+AjoH1WJIrW61DU2Q2TMgAPiz7NjyaRjU+
n83G+ZILh3ULWL8f9PXnBDdfBt2gjjbIGzz4nkKptTHxtvRtR6OyovMvw0hEnmsS
h+VWNqAC5A536MGaD4OYq3ajXCrGHYg0bDcHVPc456SStX4JB3BKrmcrvd2AgBvy
+EIET9UGxQzqi77xmRMGNvKFWSl4j/OQUKiv4PI7x+0F0kxaw0k5FIavVw82PV+h
JKmzlg18EsiAS8JvW1sI6pjEAo+Y3Se5lVC+JwtnD2XgG/k8v3yptVLzJY/Sf7Fe
wqznoLKQN/JyOfsxDWl+E6Ji7TF2QEK77DoT/NEuDmrdO8XjvQEFdDx1StoJIUTc
7/aE00r81mXgHvQsuA8VnCI2pl60XqIbpfIDjPjEMB/f2GFoUqA06y1ZaQHwDJD1
1HxC4HK+5zmyFbQK0tLCo0f89gvJtEJyIsvOFKp83LkMpMDy2ZS7S84GYqKQ1P2b
XNVif8UlEIY3/ljRJZz2+Yn97TpxOH14V+yUzxy1SyPeLvzH/ZfCDYqSWkzzXpid
KyVMlAPmHPlXV171iuAD/VYebczh0PaxYpsiqiXNovW8ldkEamg/4yMj3Xnm/tZO
ibl32R0pHszbTugFjl1n2MgBnoDDiLoMtjBP4ddv4cl6ge8B+5KmvEtC7Js0kVl0
JffSvVgvsGDP/d3TRF+zPojjqjiAi3KgRMW4mXMY6ZzePpT1yJ7BQSWJAw+lPa7V
ShFNVcsZxcvP2RJNZm7eSHIN53RzzfkCoZvxSTCBcSz7dasquxobw7yt7FCZLW7N
9NWXmtwigWRZ/zqaZO9r31h2/Z1BEzPUjUGE6J5KbZIor3wBIOTl7EgTH8PWxd18
TG9WATAGRWB9xOOm6X5JMT7JjXNcvPMTCQtkFmhVSp2kXu4j9en8jmyIbD5S2DTt
W8yT21KSbFTaJF1ULrl+D2WYiK7YyfN8AAgwjRvrLgZ72WOwRJy2hhvDCM6e9ZnX
gyvpoIRKJay+C3cHpP8qHxoxePtOkvFrCMhCzcen7Vi6COq9NiW9LKm6hPrdwM8v
LwcoXJ85EcN9hIW0rCZ+p+DP2tqNlpnrkdpDq7hfZFo8tVIsl3sqp8D07UnTFLRA
FqEDt1TdmYTOcNBid4t9W8njp8jX4PDT3MgFGLEM93cuHTPtc7S+5VvDmPCJcgF+
aHnikyKePYRERc/6wIRz5Y/uzQ6CrWCgfZDj+JMOCE1ATaPER6zhyNY6LLl95AHY
xGrzGJMPJ00CFxnPwxF/QDZHIPIqmA473ruZRjvi0HQ8xnyzgKlimpjZp3hMwuLp
ccUO3qNftDRrAOByo4cvUTcxmax6EsRzgAdPLd6RCz1ZLGPgJGdCfIEA+jjQVcrA
pQWAhjPwC8C8A4r639vGmCctc8I+YgLOD3UJSAcLsUohojK51RK4c9ZGFHpcGN73
A0YGYDMjf4WASqPTJDP2yA4hGmGzWeZZWHKrKrMXDYQH7jds9eY2wWn95a9S2xtO
GalXbETuTI65x9zNkaIGwVv9eyNSD6Whvy3pZa2pbHh8MBTPoSi2mSambGfWP7MT
DkjqLXTnxFs3HVQr5kz2Bv9+ULXt7bibfM0sLwzfjam/T3hqAyoJ1PHlHIKtDhkO
B7e78lw5OM9uDonU0dtV409tDzVyvfcfV9KYY1pZgPOAjzuLL+SP5p7HI2Qe81T7
+zz6q6eKewiPe9MZCixmurXUNQGDGTB/04FGO/i7AC4asVDNGq6/wRRTvtU7F7rt
8cJw9B0c/Nmb4GBASYoYF9F51Q42T/IPgAiH1llFoZaPX4eVH2PrG22ndSKPQn/x
BGXpC+8o82lAUjMuBBDhKvVg5Jye+gewhD/wMrI83JhvhuP1zi2QQDuXCwNg416e
3CcEiA4qIZmUxR0TTdZEJ/DA/KcralKTOoKfhR12Pgoiuz3g6PBg3VEB4lfHAFqV
xDUx3UNhZlm2HDtSk7t3FuN2PSQoCYN+7WsLNnoIlgCGJJNHNLhtgJq2E4VjqX4H
z/fgNQyVMqVmLV3Y07j6MeOuguxdoaq6vkMmElevu+4yJFLJJedSLKblXxFTHudb
aVdFhaZrUym9Eq0ZUmfGKnvMhL3iVkbAHN+cR5c3j6U0vS1VwChaR0QmZkt8He9N
MMiLJd3mhXVSUMtGYLzO7toUo5zQlXDz4zmTd+3VWrCOG9jTvyqIKzqkSDKfa1/N
5OZDvtKyRNVcVyO1DPx1VasCkm8EEgXJmovQ5zPkWNeTxUwmUjl+OCmx7KDEjOGC
EpDtWvuKnmfECTPSeUUCvNC4Q7+vnF9j4TDHf2G3tj3fSjFQasTjAp9yKDUxUcq5
CoiRwXu3fauZEfn18eLC/D0KX8ilgs5GwFh6axaGqq1nRnGjDORHn3eToN/kqxak
9Wlz95paWpHbm0nwlKrQBb9u7AxeVTrHxQqytcoQ0sVdMBpRgFqLSYSV3dwmaswr
FEW0Vagm16LA6yGX9SfU5Un2eJX7q8O5YcHYJ/vhpR48cycGKmuC1LCXEfeuRZTX
PdSnEkpJt59/91TrrwPSGYC7I1iBMhkvsxcOA/E9fHRpp0DUTF/fKtu0XutkdoER
yQWxIejJhDg+Y4FA36rTaAiDPvL85AAjn4oQ5eXPS0/dwvoqPLY27m9ArxN5EU9o
rdmNSb92DdAgin9MGUaruRL4kfKd1x9lmr2EyVfuIUQYWcHwEyBqr97qp2WiOLyI
U/pGckju0L7s3FK0PI4Jw1+3AZtoETQwaZGI5vwzyv7vDe/9gNUtv/wGaW5KFsfo
2IZp7e207kOA0TzLOitKE9xiE7BVZFAmyDuwvwpf0heA+ioBzCfDSdUBSn1WQFiK
ImH96QAXOmN+XeUA0/BS684h5ARxSifcSK/+JLQpPSSQzld57VOx+lc7ztQlrD52
R/HNcRo5uCqBUUai+Dls2bNo1MJhDQcfqGnWBOlRhKEdPbzEtr2MO9xnknhrX4CF
WcZDN83C0I8bLbwK5h0qPnUsXkKKNOKAa6dHqiM/SkR8HMp5iEs3N0JA20jJn/zi
Xguj5DPdFo0CAefwO6b8EhNdoZEzEjCSzrBEE+jQMtHHLWE/WTUCymxGhC30vmYB
gyJ8TnbHjxK9ML+byQZm+feQrxE+NZJ15vMwC0B+jE0N8hT9DZtinL/LKuGAhZir
mUD20LF1aDcY87Emb+M+sbRfiEfrgaGYFW0879DUNIo1XCZ/wIJTkNFogMqXTFvu
O9evP1zEso33LVoCacosP75w1RlL9SeomlM2ZNNNXTVjreodFVHtGUOvWXqbH2gO
uwWMVtDVCa7+v6skiCEDFRK9Lc3ddYCy0rhm7RWtCnzv1fYovniWsW2KTE8sXwY4
mY7NEoO0JOFbjZdYWqAEG3hHFhNRGn9/JhEvfYunud3EZsVRqDwYkRE9NEZPyiHU
vn/skK0LHfPBDOoJ0nu5d/0NOpmPjJEbgexcuMWtHddiPcvsJoQAZ+IoEc+nbXrv
34fhOnijxHA8DlNHg65OxwV3S+NSOd/RQb3L3jJj/cbfusKBUub4j4xvtRx1i7Ko
5dqhLoy71HZ1ij1PpKJpXhd0vdSjVhscaXuzanT52FSiZGChdu5Ec5D1JynWV9/8
rHUfcchDYfq3utNyvrQg4qXg+ohl6sVkZ2yCNFaghZSixKI+1v6Ej8P2Etd2ICZW
VEbLWxy/B2cMeOxUebSknsYs9SzkxllAgjEofThPVo8vOlk8JiXtbIhspotFg1eJ
/4vcNnl8QKNETxn0XuK5rouN3UTj6T1fhZK+lW1AUud7//GVSFPUXeLQLmVC9rno
oyZVBtJLA1Kgem68k9Rrk89/Ah/HNOqI3wkpZtq6CeBV48bdCfw7vEQY9YcJ1iJ0
zu0D8uMqnqbm3pBkv4h5+TYVvK/7oud4CpgDT+WAAcbw/UJz39l3w8kyFSH1IMMW
vOrzc6Z9fq6OrMKd/AqvICdRgugRfvRpY7cz4wfAEGWFmfhVPD4DjM3/jPCD9+Ov
I7ZBiLXYZxFntw5E6eH4HGh6Ib3bGvulRHyXVjr9HaOBTiuINpULUlyp2tkeugaF
mFf1ThiJ1CjHXjBKfZR003SBQX8QtMGspDAvEef4VdhtrmCvh/VmFsIhidTkXdDM
RtbzVJh6BUzXWWSArHXch05yUELJIJKNm+uZmqdlG21XUKO3qX6F9NCVkXPB8duV
5NVXY7b2lLVcU5YeYphupuXhy/4ZIBBIMM4l476lnaGHmO5rahqAI8cP2qzx1ykG
L0nsDvlj63MRiz9ReP4RmykeTJyr/Xk7BQlYptJ8pV2px4RSE9XDiQtFkszDJFRu
trBLsxfleh2YJKRFDb6C5g5SIi8JrJcYan+o7OnkjwwoSw3oXYTVB/ucoxlUkoFr
QvgCdqDvj/JCxVzWqOmcxKB8gFT6KSF1JzCftoEzDezmhPQGypQ6NF5yKglbr/TO
tMVHtMcdjaKQ6JnLYJakxlOzZ0EwtqKRGFrLWD7d+ZUe9NgNZqincVrlSVJeNug9
+iq7t+/7yoyYrz/mcu83n7/o95f0WUs53LQ4yigPagcuDDPCzrm2wYPbtahtp3z7
ITnRVSs3+hFvSZDTjjPsdocwn7d6nDTEOzeB37FHAN2SqC+elK/9u/PUjPp+3KVp
o6HOZ7vnZ/ARHZhqSixbmQ2FP1/jR9skqyzFoA6n/uN73wOz2iHLjdmJ5GhO8vOs
td87tFaALnnJyOMMdvYiUXANkyooT6FNZ61iGajDrO8HqnA/64Xu8j83fEq4kVSV
gEMOJOyIjDFm4YG2gHxxCyc51vOa86V+OqZ4uLeaufSEDYkhHbdHu2qk2XDVrfKQ
0rT6a5l8q5UmRs5ooUbBJCamjTIZFasAczj2XJ2B44pXEn71tWBig19Wb2tiGECB
+aJIn3HJn0/DhCMZKZJQ7+dq6C8ER23eN6FnITqpefoK7JiXFGbM82CooENSzRJb
88tgc90o7ceUAqdquGcoo2qMsLMRQsaIQDM318wa7GCQI5KTDPCoxMs+X9XAyJR0
DFRzcC/NQp70jGuIETDQiBTtw7as0kBuhY2TQOwFfoKaadtwJqKrs83YNyAdGq7F
86U8cg4sAOqd0xWprHciwmoruy2IFxc1kWtfqoARAvnjLzY4SaQBbSlCEHnDQkHw
lX94rc2HgsRfmTeDy2kY0TUSLZ29lxOAKnmpPBWkVt6k+Kmnbh3yIeCv2lgjVT61
icnR/Ugwn3pnPXqc1ALe9PUDvHVQgN64dSj2V8iGaHSI48KRoSaft9WDRJS+4RkV
8xwnY1RElOMj1KXpBEx7UGyM0bRe8SPobrv1LRhe8jwWhT6nwNXEJy+Jk2MDq9MI
lxbWknPLI7/CotOiPvfpbzIj/EmAvo05f7UsZ0SWUrzZs8JBYpulN+OqMK+tbT/Y
obFING4+jqdhj9DIEofH8oYODq0ltEjOAUxmjEFj9mq5Q86BiQqlpMTh0A5yeepQ
cMujxeN47LzIYrr2kXJpfQfxS159Iffj416piXlxEZdpxIO4CUjtDIZBVgyJP50Z
UMqTwo3lV88pA25nB3ipCyWsU65y2/JY+A6QZscs4h54pCBeb9g4Ysl0nz2uePWq
MJE6YxCHgIdyva17Th0tGmgnjpjKtp6OJ3S+PxNtJQeIVjWQxmDGMhlszSwY0s5x
uCgJNi4RUia2KUBikHB9Kvl+3nT7s71FxXqk8g8VITxsdTamh5eZOHrozQn6leN7
tuLWzyPvNfAKXdzKgDjk8XFVA/3ktmf6XNeMz8eXbTbCayJwFMdPXy/HS8KeVNwo
7UH2fFKTtY6xIELkKtJ8e+pxHIOCRmbwSwtJMCpGFLViTgKHvnYFDCMEf49CmeL4
/Nln8AFsgJAx3Zfmx9TBXH3vHASBMf5b1T6JJaXi2EKEwIXC3fk/TsPikIVD7HgU
ye2qQ3ebnZ1Uuu594v7OBS2T0dULTyrtTcZsdZCyfabv0kLxsWPOqXwvO5kjhRvg
6y1iotOWFPK5zJtI0U7nMpm+WBfx7eVk6fyAQKBXE0kpTQ6Y7+v/2a//zcEKoaoP
y/VF1wm5Qhq/+vj01/k/0t8S8KUnRwhnmbh0EiKo8fsTN+ZAwa6iXdMltN1XbtuI
bhoj5s89F4pDZ6Ij/po9r443nweZS/k0FajGcumEEoue69PwKWon9/aVOLqC+pQy
/PVvybkOXmaXZC71WOMDJhd3xvBKW48aceMnnUtoBlSkJ3hNZXHMOEazaVDifxpT
WnFjPegKYBYB9bxaV1Uk62h3Z0k36VACZ2oi1PoSLvt8KxXtWTWP62yq84/3hgY0
H058cxiL8R2ktIj7lvvsdbGWe6Zbknx8VB/906ZdATSFlDXrwlUU9CahsQ4A/ZTW
X4wCa+xnwcGYGSZY2d8vrgJj56Ad5AjL23Z3uKPZmExltqxtOWteeRZkWGuSpkP/
GKi6a3/Qg20gImiXor9HwNCm7PfmUlMRrrTJPAwnv4jSjUhbut1CfbMzftgAK8tQ
KFvImMAsnU2pDXILenJY7RFwarIQ8C30phaYksCMbVwIJ0bIVU9kWcSbOIi3t1dU
/kFzBwWiqD7n3mfI26/bRABhAlhRdaAVGA1OdP/SkpScCcYeo7FcuIqYqEG7TvF1
F6I25bA/xWJUHULgk+7xtvpFUl63Nl52CyeDavriIhfh9IHrxBfXU2A53FyaQ4tX
3X2+QZJWZ1oNiPVfICFQ+d4YgKYr4G+sfQFfn/UkV+yZCIVQjvk/hBJckoqO4ffx
2NfFYtDk2gGq5cX0j7w1SX1Gt/6WhtptV4QJO8TZxyow+K9H0OyLaBZOyQy9W6YH
QnJC+QfiJzIC+1WTbqPpBkeWwGQfblhc6MKjWVRH6xAbNJW4+e0ehHd7ORLcNq5+
c3MO6qRb2efNRNkVDq81uqNl5dBljSNSwAE9xSPQG7wbtAAJ7D1K7yAJWSwit0fh
krdIYzkm4tWakh2/PUQwX2wvC2TmRx0BDmBNO5liRMqbHsOAeSE+ppqE+zicSyg1
QKPDyckQN7twVNTlM9HvY4vQymny6lkaRSQ3sfkjVvGjqOunUF1eZOdhXUmID2fk
dtTMRfr2vtrVGw4iHvGLeOgTEssfb9C5ImfBf1Y7i4AvlhsQpQMaLQ3OA1QrmFRd
mlfHyugrPyydaFZEGP4qIBvfEH3q50hsH5FLf9q4TSd1NCTgeebQRsGfmsEZzs/5
9nYmFz4psv9W3yXH0KhemmjLhkHrWmIotC2bpzHtk4zctNv/RQzeefwwuuD0rYW/
5zybOoTH4YZmORAdLoztS6JGiTRFrN9U+2ibmeGbTvQOmLBBNCyt2Kg/h9h3BEut
nPK0J0YKX8ekclBYHsxgB8mPW33Yau+wXcgR/6hMjw16SXl9kQSLS+T7pElXZSlJ
yFcp+9GRYmzQXm1zdpojbP8xGc+WAEv2PQ1hbzrRKBjqtvxccx4V3XYFSucAsgHJ
Aec4eMF8j0B/e1i45TqIcm2VImRu00ApgXvZz8e8DRfCuPv16Eo+E7YO47yBFKoh
datP0mAVy2JTCmxPWUbzvn4vX/uGrstIoMNI23VECUN4r03lu0AtnfDYyygMqWpJ
Zim3YxdDLWh4QhO/znMJJKdp2qzWy7MjXfQ+c7NDVj/iM3hzcFmkKA4VTZ29yCSr
u5jGSTgRhENC0ly72IBUC+q0x8MWaBpoKb6bNOl8LHOlCkxPRb24MDAl9iAGVdGv
pixZ2muJ7MzSQe8eU0XxxoCYrlGl5JhEkIN0if6pmqY+U7YbiEYt3QaSgKRzyiTT
amdjEhb1Qgdtrp1sWKSei/GR/5XNxWkbwgk97qSg2EmMq0h2z16x9Scbc67qat4g
2NvxItmqHMPP5m0mM758/TKLAGXMGKfdsuc66WkzIuN0vYdjOcxgrLwH0Uw6BjYA
MkUH60UAdg0AucIrnvieaP4uxAO7lZmDMu9rG1DmpEfBGK7LaFDLOToLYd80aR6P
Uu8ppUZ/wIj624YNZ1qQxDFTiwizhep8xJeVJVYDIfHUr72VCkG089WMmJ27H0cx
zatJCzmWy/oNoCs8XiaXrEiqn+o9N9YB/BXalkeavRDHTNzc0rqm32QGi8hdePkI
uwQs6gzlTKqsp+3sAv/qpudd0+PZHdsfOjeZrj8e24bLsZtrZOn0pNA4s1eIcfaX
FMPaWNgtXabuTw4wvYKK4ZwbcpRUUuAmJuIRfuAbYAg1W87ZafRHO/DOv/47S/SM
sSbKCNV4ZU5zbCiXt68ONMAxKwLyPIk5o5Wg897HSOZKoSLHzF307zZ7l9qnL+sA
fbeRexNTebXsoUT62zWIftYUV8kCzB+IMoxk4CR8anwRuHO5xC4TdQJHLUN+B6bt
yEjAQ5DjmN8vyIfxKfntrAzY4PzxvL1B052MNQOuikNFacvAAxj8ess5/sXhzaEA
O/mfsTnVrEmmXZPLsgD1xr7aN+grT2aPWxk/crsCYA/ucXIVH3exPWE6F49ji05B
QzYdM8inpN6j7UAz9gggUnfZlegmWR3gT46pzCDK/Lfxv+AgojuRUIcHN+EMkIdu
tG3pTGlzlO3+G+RKFFQ2ropYUHanuFz4pJLUM6p2M3NV2jevmF7I94I72yG6PoZa
HwbAWBfEGJ1TgzNGXtK9eH43H1cI/t4rfV8bk23nqncGc2NBYDz+Edr1yBb54p0Y
dSL7IpyM4m/7UdN8cXKTTsn7TWJWtZsKOP6D2pXQUtUQVjksfpyB+N/yUeu3DCG+
HS2O7ZlTzVdJik3eZukoF874KP4itK4oRLZ7c6OCJGdUJ9EM5wmyJ62bQKriUdSi
eJAe7UcAR46MyVt5U6MXUoMF1OHpfnevcMyDuYa+XKyN/WYK9kZErDCLuBY+Q7Xf
aBaiGYBmUjHTMVJfLxIJkUx2k5SKNNtPiQntr6ZJEYPgTVUFbis+LUw0VoiWAzGV
10F/ye+yMrjjIJd8STs9T2fk4YkA/wCLwmX+7yr4XgZKraP48zdA0i7DuebA4e2H
P0FkWyQu9XX0naZJYTK0xgvz7L+oOJ7Wrpqn7MqryPqccnR3sbkEdyK2ARRE4upN
ta5uOKei24YqTnzgDd4XTCophOKXdc217PP8xU1+lH8u2mPcbk5QHd6NpTG4zXzc
3sXVNYyrdq/dp837qz9sUMUJgG7lqXzzlOocrhSgBtrRDSelM/BlWOB/CZYjP/AD
c31FCluZdcHrTtXLFu0o3lXiNyBKy3k3w3FNCRwgMpl6KSy+m0gQ7Cq9q9GbkIpR
XIZ3YAoPGVs5vztVQ0AI7f7bKPGXAj+cG8Hqvq0TQ6NhavbWqqAoJ8/6C69Z+2/a
JcrSfquyHd6wmSQMScAdoWtZbm3asiyqx+bRONZVOeJH3cM6pcqislLm7vIKAkIz
HS9rmA4HXyQ/AfQIc9qaKK3/LyMMuxClUopRppHz9LrHDLiDazELxPzlK85XkIfu
qYWbUrPlTlcNZfRpPsLKIUv2s5KOqI+LRppYiuy5siZIhV2hPSND37hsVo0fQuDD
q9fgJIJ2IHbBFNLdsHtQPzabGfik9B7Dn9rm+9XnAss0Su+fUYN/lkWZzTtBszNI
u23e18ceoOisoMI+TiSRkm+FXag9LZj3QJl3x9yCrj7wixhggHmspj4tDEjAAkFF
cccggVzpSkG/4v0MZNPXw/MrfJyB35x2WLlyUd0sSxzDZ++SepiCBZuMnWLZhFpe
/x+YqPlWfatVBLTkP9wP8wA0I3vKfOQ3JSTIYUYEwtoDKGxCOX+GNzUcLfWVg1+l
EPHLk6VtuVpGqTlxPrEwGm3Y7EVH7atSLAZRkn5RffxIBPP6Lj4ex/1Qkno6oMGx
/kfYR8mFQr6+4FUvenRtZNzZ5+z8WSvKJqqEybm+GVjlvglfjs+YKbfejW1lTZgd
0L5by4rYwtWFtLAAWoyau/iZc7Y0ujykDAS+1YzdoewREZ31u5ghKE8/JNOqjpCO
S9VTSE5aYLCPJAu/1Oa7P6OkYSEr1RF0FrMHWa4YaCA0Hdx9LQV9L+t0H0thfEsw
DxRVTTrKbu+2E9ps4VxiMsBRBhggZuz0pIrVLed/bPDSWry6CepVjxUWiREiIVhe
c0h7jmHSRR/RQIH5YEDGCqmC7SMctoMW0nsUcpQbbuyhyXWVy7F5h5/PKGrLGRcN
f5Nvo6oy3VYJQAlva1q7zqBWgwrh17/OYkUPc9Opy/pJ4LWhR2MnrqtKXAKX8J8z
YRdTIK9RAFNqCwDAmkJkrmm/XvMMxcpD8X7YyWrWP20YYbSREZHorfikPUMbV03h
IXqqLDWhL6n4boH/RerZ0ZjcVo/nRczVbBqYiGlFPv5YrVg2+ab/vC8M9XwPx31S
UQmYMzfqZh+RxCRiXALTLfE1GS4UxiKqaq6lcNtEIdfEhDFMT4f/9n76aOU/Ccmm
eTvJ0iE0G4cgS1tzTHDxPbPTj8eaMkzi2aAL97I3ZKmG2VGV6B0Re9X/NwOfcYkj
v47i8+YVs6thmPgAGUw12gbJ1PcVi0xw18wM/f0nGUQJwerTQZmRmSyxHxEjoS6A
cDJ+PS0fElZuKBA5O1QYK4RlK8OprsNcVdWAIxF7X0qx7O7kZYpZtrV5/5lWtwJE
HNz/p2zyyu/a/owF9hAANvZSrNHvbuMqGURTg6kjFl+JK9RcR+GBQDo1pnSnfAl2
iX6Jufc3XVecgzE0ca0jbtXllJQdKHti3yf6Ser5aW/V9kapxF1rZO4Q0puyuysm
btqxXRIcBwqaE1eeYySmb6zDbuSn/NClxI+HYq2baP/I8qczQagvsc1zFnqroOkO
ZbQTpfE6o+qwk8DwuJigJAvVtOJoQpqgdewGBk/ZRZTK2+ob4vmOyd9LD6d54KON
EqBHb12H3EtPGx6EcBskItfjV7ZBlctOhITM7M8y4zMHPLfQj4GV3ex0C6+TfMfA
M1WID+nXt1RwGLXH1v6uCdRonOcYavdsGtgI6AqiZmnxOVyBzIghlZOjmd1X6Yis
4U9WJLXgR91YK8NmozSIFDGPEFUWm5Q/0cQDAsi1aMHeJ388SnHZ0hjsNW1RssFl
ZXrosT/SKDdJ3NXHLWOQEIZFHoqX6pnE/ZdQzMJuccMP97gSwizeEifUSF58+kVh
mPhtCn44Sfj9GV9Is1x6oyqwkdmro8lba8QZ2JJHUzX8rDmJk9O+g0oPrzbSuMqv
HeXYDJNUikIqT3xTQgKeYzSRucr98k4Cpo2dGPS22hZMV6vze3ZPq/2PieuHNpDO
DTZ5FLpRymRtQNGczZ1EorvGdJewzI4gmJre4sTqddhfoaCbgi0wBUhPEMZWpl+P
ya4gnXLpHdrwPLAq5f6MaZ38yEIkrXI1hW+3bGFH0+W7SpKDS9kVYG2adfNfXaug
C779MgFCTW0txymAZNFV3zIaa6hULCebvTf3KZcrnytHvzjpJU8/s2ciQXKbYGh2
DwATrEYd1ja1TBfNfm4eLtLkDHX4N9x6rxEKozfaGXq9qw31ifrbWP99zrU7wqQT
5bj8hd2px6UiLMub5rs3xk3yLrlfovIvRwtGZ+8dLVv4NPYtbz9jZSGcYZlh9qOk
thL1PBU85MJB1fjeSJjmtngpPuHdLIhhwTD/6PFpz6hC1kdtME3FVB4EQUnI4EjN
jKWOWMbToYPvsHCdOXQt1LWAE9xF5dRxhkt2Co5HBPPUOjr+4ZdBRMC9NyXbmOQs
hyALkUccdVRrDGr9hjrHVAd9KvuMd4p2naOLi0+awDfPLVqUcIZtRX7BTU8RcP+c
1FOId/l6mH1e+0tX/C6pKRVaFJQqA1FbU4I+hfYW0r6p3KzbMBIZij4DQ/48yzS1
3WHAIu/QY7bXe0fV/wM4eYUnj6lHVsmF27PThoanEjLbIgBDwLeAQHWmZf1VIWUD
47fiQaDEhvd3QYQN/uiFyJ/RoZ8lS/TjSbjfy5dFIpohOaVI4ey5hc3ziAk3iL8B
NS6HM7YnARJjf7n+DSoXR8y9R2iKvySjD0Obwo18kFK9jboBdSO4LRhTGbJt3p3L
op+27NPq/hvRI12pkdrNx8LAPHszFRIpHFEpmH9CPYRgttSGmECaAGUMYCCFWpY/
JqFmKZWQWtKTsPqFyO17S157gWP9iMbPPIg2FoctvtZNfF8dDj74XfLQ2nEVsO/m
maKsUi5TXP29Qq9wrqcybe+xk9Cmgsc4X+s5lVBwNRnZGOL7XfJOLpb41yceWAkD
Um4Oc0wwJwpzmpAwwdd3dVp0tErLew8YS7+lW5h8hdyE1+nMCeOmtOm7tDFOtzN6
roUo9Y+UjO6MjHv6ikv4cdFDIn0otSjpa1x+kDnQbhCoVFn71ssOy9gogcOKPjjn
iK9U75Coa1qiVhdPHDOOGIVC25DxRwiiceU423Q7S8AFN9Qzno7e7wApkvfW8fBX
It4hq8QncElNZLCalut7IqZ6CaMoRPmulLd/rwgAFbkx9i5oPMgTL1WwDZfqwDH6
yda1u8hXNfIqa7oTiohloBc/zNsTtaR8wJB4kWwqa1TvJ2mTBNb/KyzC37ihSk9b
S1IXecM8RTHmyBYMarCO2R1n+LRyhm8Daiz6EEB9d5Sew+Ezdsry2k5zjgnT1ZCV
qdQI2Me7oHKH+W2x29i5Wd9kMuO4ItgI+gUlM9ea8snZ0k4kyHzyJFZy4w9rpEfH
VFaJM1bqBOetROABxAEMDS+vdx26jCRcFT54bKM4TtQOXGFu+NQIA2zu8nEZnm74
Vo+meh4DBENJr3hlkNnIzQT7CkCxcNHE5h/wr2J0k6vu82XJiU7E0fTKE/uAIFWa
m1QVv69OnRHfkUX0baT7uYe0I36ruIaNv5GY4lFylzIgeiG426tOX3+Pbn0w5fyl
bOSbFrAMpm9QWmINPorbiXIy+JYKXe6q8RBgdAUgcmr85tzqM9ZYa7RfyFU020OZ
MJvTJSLAqgF8xXtd64Tk8rMzUCbjk+10dHZCeEYuw5GgZGaY6Fq17oTLd/vUANGY
GXSve7C+AQo66W+lJnzYgmTAZ8TVfeoMZCdVka0SMxw1Y7humLA8/zJ8HKhzUkt2
fmLLoUeTryA3sA1Qi/5KduASwOJ0Vf66gCEHxr2H1dxWN8w0tFiL3q2thK1JriEk
QVIONxb2QJVl0tPZ+I/7gXqvx0vznTXah5Oqs3N/WyC1pMvj+cMeWovO5KI8aBsW
Ec5tQQks5SaibcdHjmLxKp8oDJDp4DGCrvSG6tLCGYxrOHincKhoX1Ebo53dmNmI
bQBqx1wY3EirNXLU8coLtqKhsWz+p5ODvIMBxptA2D0CKmFp1jJ9TPaP+jX4cgjD
mmYJumk5k1R3+5JkkNU3xfeJwzWgpm4oWx5XYNvX6i0mKG/IriqoD55igbSvHkRD
My6r/8FKWowRyqrgGfP+OGvfjR45Qm1I2RyoPoi1MVRTKCsjs0uAZ7TKfJH+1g1z
pkth+ThJty/j1bhXMUXr1S3ZdWHubm9rQceKElTrwgwEcplkBE2FFG9tYPaEjfX/
2eoMIsue54/ka05Hckb+nAeWD1f7+Moh7lCowijU7gyYFTKjqkH+23iPg/we1dKw
jpOYtwW9UxjbqSGcmRX4kZ9gViGKFBGeXMXcUB3lr8qW/1jbS2gaQEIiUJ6+GfXA
MPZpkKkm1yzTnaXJmL5Xb/q4blA3MP+gkAKhQfYrB4ZBaU6r4FxTFnk8WSlWoQrW
2YCBjZaoakFvtP58+28GGPEwoT6T0OSyB5VqVgETnImbY7oeGXhDFlx+8SycHwHr
UFJA+OmPYlOQ+aYDbDU0Z61Yuon8L1rB2FI6lI7riJULxPREwpH/PcT20SxDrQ/2
ssNP0cTzf1BmAW5cLennK9uvPjhm6u80i25AKdTDX2ysJU7UY2vNHkxGWIJvI4Bq
ru+fSCSPiZ1kQIBf3ZN8/ZHn/H4K6fTlpPLPnfXOJIRYCzrjCKNK7yAROqozxuXI
2PAiu1qpb+gx04QlIHgKdw0KoORRFHwsTeDv1PBoje+mWTYVB0fbmgacvElVaRLE
In6WTlcPWzsEtkSxUIshPfqH8NEvVBAErMeK1AbBPAN81284gsx+F6m5flxpMML/
pKCdrScScKGGXoJNxtpkZga7CMALbJseJOBao7O+Z80/42aVgl4/ST/JGBSr5hAc
LaS8nYM5FiVSb/CE3/YMC2B4UCHRMzhumqm6IVFuVXhx4UA6YG6uGdYHUYQr8mQK
EcjD30xreg1/Ek69otypt1mC0uEVjGnxXaeBcUcjLgBggsjYAl6jz/m+TXbdq69U
cNsIG29L9MA3n0qs0bDSP0fyqm+p4ImFEUFse1/2PxAV8So4uWAoeU9IA9vXOX3s
/V1uj5CEpAyRdF2W+jznjRhWbr9rvoxUlGFM/b5W+n2nCuLHaTsryRV3Y5e/OVDD
4GfWl96lsEYjQk9w83zIWTdWspOEGG7++0JCLt0aBz0LNhPiZO0Rumlas9fFq3oM
lROT3HFjMmiKlxhXznKd85IZpw4R3y2LHu1nt10mxQ4CXqWjlMV2eLpU7H08bJuc
r581VNa+i1UarcabulGZ3ngv3fH2V9GmNllf/UqcaLgF43X49KYdaYw3Le8oIlkG
r6BJix/IeMM2MyzCCIj4PvePBx/a4Ac5RcHXw3cy+RsZ2PPd5lbh2n1i7QmqPjUG
U2uOPiMvEOmCzSxTNM/Gvup+/dsRSMWiX4o3mYXteG3x0ypEvSRDiGBz+9kU22bJ
Ede5+bnStwjSHPrV86yIBbpmH0vajjVIDo72Pn6n9fe/BdUiWwzkGsQEhschzepm
E2oRga/B/kun20RGLkuKqexyMRJnjR4lm7qSZRpcW18TywAozV49T2EW2+S0pxzj
2jpoOUMSjnNJSxy0El1IFwafikU/yk2OWMUXuok1+/J18Iv+L4kKM595qqmAQXfX
WTqshoCsqkUhVajGF01qRZ+Sc5Eao5Nys/WM6tpgSsCPLelngZqNmh6B0t01dJ14
WH7KjLQEtSH1aAhzTFrTvdvJ7hvdkkDKJSAy66K5GY+whxTqqI+/5R0SD4ZVEigl
w4aQKERxM5X2N66GcDQMKxgfr4hgGUUz6zsfa44Am3dEeHCHCGmvRT/Twl3YA2j7
5zLKAmljFji1F3BRkzIlWjl2UysBf2fKKMEgd93BXnWnGvT+3jDKCc9bVFevHc9j
CUbMdRU2Xqx4HcQWgY70QB65WVspNJR4Ka/+58na+0ZwcQ5g59uN3fC/efx5J6x3
r5CiiQHh8fIu75l17FbiZCpP0G5gRbuCgVvxIZOINzNtD54bVRs2qj1O6YC7I6AZ
ZA5EMf6Op+wR23owuBZfam+AAMDJUpcglOz0t2ycsGB16a3kF+GFiz8Mh4ZyF0Lp
NEgdK3jZZixdZlF5EwVn23Mk3D7TBr0hmSKhFBLWDOJ7kzPP1J2OsmB7yio2RSZW
Upg1Mi/+9gFcy/QI6AFxaPcIHbZ1+5jvBQYm8964ujgrwGJAcsV+wewf4uwwt5lT
9/8/xV1U7uSaOXckB7BIlsYGVObqqCXPDWJcnAZyv6fe8XHrc9lFdXpHMO/AmJAt
Mgxz2Kqcdts8+zBZXiRT/Hl7RB7v6FkG3aRJRGV4sKBXFaGQrZ09wB5D3Ia7sraY
gXV55FYw4ImNoSnW3xBMzLHPb4C3Pn+zTFfMT7iEuDsHb+kYI4cSxlaU7M1UauP1
OaE/nquFP3h10up7OT+Ft+0lXB6cKZg6uI86qFtpTzHDhW7V7Wm/kxrEtBY0xqFW
hBRwdV+W/1iNBmZYwqviIEoEMRIVPFUE7P1TAffs+OLdvJCQIbsMARjxXugv4C3p
5/th3E1LWxqjxk2UxdLMVmvAVXTAH4JhELU7qX1i5TQFDQYYbbE0OjD1q0B4xn6P
6aG1aP3YH6T//HovwiEPu/rH10GsZSJCfmpMevj7KeCwUwGPnj2D+DDrm+5o6rbC
3rWhgMsmygmB+8leaQWMg6vSwyKc37tT8DAmwKl1/k8KsIxfTw3xUc0MgO5MitJp
DXc48/r9RuVfEPFL8Kv2nCu6PAIJTnW5aCFQMm221DRmdYIXmTM4I2xOTqEe2qHf
NcIIpflv9KVpTABaeonbB8v7s/9rIDDph90GtoGb1FIAbw4xvF/QOo116cD/tLv0
gXt99nes7/LiN40kFVxjakU6ps5qLWsmhNNwUi/QnNBOpaYSZkLzQMyUZvy1vCNl
4CmQwKJIyrrVTxOv74s5h4DzVFbHHfI50g2SX38eSwoOHJIWSRTid9jUmhos9sMy
QKcCDUp3n1K+swpcSaX5Ri26xzNbQtd7hK4/fqmIELOLow+ORnePR82YoTWMdSnP
hEQ2mQDJ6+jLXzvPZUfFIKlJsaQ90TsXotAtSeemIz13qg9A1zTAAHtex9Icva9h
`pragma protect end_protected
