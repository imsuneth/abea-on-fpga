// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:46 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nZNOphslBUnosuWOhVZzI70gYcg+oQfsSXOgaTFzpOwIExUuMxfIpRY72gX7WV3L
BCXgXGiss2sOljKrFy9JKzhXEiCRRFOcebcJgBY18v93xOYjjXH8jkrP2t4qfSuz
ifH0/EftbT3JNyQ4IvUkqKAyDzZCnKtb0PPnbDwI8CQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10464)
38aZlEoaB1RasPVKlU4rYFR6d+zrGE8JrEod6NC5GCG07fYpiqcQM5v8mnhtp6hJ
+Oz/I5OoQQHdDnXcO9S+COZ1O6E2cX+F+BSqJjaExX3DS7zNapmPL60qn9YYjJZd
q7gN0IqimEw5BBfq31krn6O5LXa2F1XThlP+oMpgnuwPMJ+XbolBqztmVMqVLsB8
BxjxPokMW8bZwfEM2HA/+zEWzegMV080mwANt6CZoJG4kmOx1ImCqf5a/JNLK/Wc
zx2uhCq2zFlH+sTjfGKuEe9eqAGqn0LMEycu54DtCaevG82VPRO1jz+75EcjMXDf
QSSrZUxijUf8wB04AC17C+WzwlykmZnYb9/O6/Hk1+QbZnmRxQXVNiZ5RWbkyDnf
aDM7OWo6S4wKC2q9X7JEl1DRnLqA0lOfXEJ69Ped2xMI0Z75wSZyO5wLUeCb7YL9
wR6oUw0nW2yGAV5Xd2W4zDJe3g1nnHqZUnvzq4TpgaxPpohOlQmHwv/+pPCvY7uT
2ZiqN+/Hv1CMvTP29iPQwsHG8iwG/HDVCMG3GYKIgtiBXgKWs+B8gsDXYRSrknZl
v5Qyyq7a8uDVBBf/foxcEoavNjztEkKEtqn2neHR97Q+PUEBcEwPJhYasyr+/OHq
IYtENNyUTIlvvVxUUk+nMBKGdN/nf5LyN70tPYRNohvIoAzDaHC1uzee84iS7U9r
M1adqm92W7sTnzDFIwRXgYZC6Nqi/88jWJ2lpIeglCT6h0pKmc/y0pwh92vzF0b/
3/EvIMsxVcnw67gDoA6/Divda1PJuVODkoGglwarkh6cPmwJ9urd7AjDipMc6/ai
nJM1Ddh5q1yJxUeqE9oglUDr9aJr/wmihRXH5AyZ/D8Zqj8nEy1OcBeXiC9gslRD
/JUyJulEhtko1uPfwHn2aY3vYjkhGRJuzIme2HcoI/h9ckWxTT/sZA3KxS+UrM+h
9kbHtotMp4sgKMDKnRCxn+/SgwubMmov2LHkqRstUSew1ze/Zy9RtidSuG4iD+Dt
XNZjh6s+lKyBvgtzejpi8DcJ5TebsWaGMJGac16G8e4YIe1iouU+syt7I8yEnhKE
9IkNQ7pN2AwVvXxipWc12mLBIAZyets7yWa62SN5Lnq1NBz06SkMdMFuGnBpDNH1
au31gHUYt58yK21mudsLkjxd0VUBoMytKQnNSwbqdN9x9ojq0gI8QPQKao0oH6Fj
hgBDJPxom7Fv+vvH7y6DSR7vEOihltz6DYn+RSE+EtGcdfXEcO2nygVpDEUlv/Li
w+JulrUXlSvNJxkVC+7g9ZgzcjNH2RVBws+LnG2iAVmNHGs5D+b7K0MiEwo8RrXX
XPh4l5OZzu9YcxDl8vIUt0DjPvdxeyVT6z6W46n8Z6pmqK9ihML2jpor/a5I4ttR
eMxW9MTIjqB0SbqdWsRiX6cNqtMIfa7Ss5lh01Usvzl5YYle2Px/5rUyANgjc8uv
DBYyxkPCl/HV8la1/c//wn+EM+J4429FigRWNmNyHiAxg9v8hgOWOS1jm3P0Jw0D
FSB/9YAACNbPyIKyVNU30KE0HMop6/eXWKbxxJt7VlKMui6HlmJ2qNIpFvAL30sd
AFC7xld43N9odUkBZvhz+aB1yeTGdzsMXtgPTqCWYhpn8DvIXK+akr8vYcSNBb+L
FcFVhsWMqvYXYemFiiYIDZP3yr7t5VqF9hBYrO4zWBPvZyW9moUnHOeiaHLwDYH9
mI4PnH+wDcFtivIZDT01mvqkllSLxp5tOG6Q//+4BlNLAGCIdmMV3fFkq82FtLVO
UzOEoRlmTV2w52WHM3+YvhAaYBBCq+z1WDiXqfv9Lsa4VsyIKqCzgcya4awrH3DX
z11dPbIeuuRumTTZdmFOAA+BhEnXDaAnj30oVdwVLkz7dvGGKjVWUA+ktPnWXugF
Pudi3ElB60ZylirEwPBkv6r8C9p7cYX1gq5OEyHt1iEfAz7cjN8vpAEnIuTfj0k7
AHrG58ubJePHzNZJF9d27H+jkQud6vJhxv83QEBUh1rgM+qXK+JaR1Oj03ljo/Vh
ooAB6oXyK1Ce8EPoBdBoiWmQsb3boG10QUHYV5MtimUeZhVQ3y+1h9MYohABKraX
NrdB9LkLVkjVvLa2sfnqCvELZ4cLpQrMnguHLAEhToOyA2OdRSQk28s4gFb4NX/3
3lfcNgb9ffmM4YRvq/YVqC36QFzhrXGyCUWrlpU9iu3a5qD9+JluNhaaXvHSOIKD
K2M8677uHCfZbaQF+r3tFx0PqNnacH3wl6H5u4feWGZnz3F1m4WS8hggvDPhlSSe
u0/vQyWFMsxM7lJ/UhtVnFm4NvBwYAxju3jlGWPvUoCMO3PvnuBaQSgR0MgVHfL2
YTFwjusZi1IIGeb0pA6Tz2O507gr5l7Lp3sM9xB6gRVRJDsLxSk7aGe480co5heb
nb3ZvPUpar3tgC3I19p3HzTgS/JJG75YmhWaBZ8QN78cfcqmvwitxjN/iamFwhRr
RWj3sSp/GBkp7ygR60FPbSTE+T3DTy7aMBwSYqkNUnQErWh5gqlawjlo6O/3oolW
y1xIEVG6JISyPTC8nFGf+cmw8TlRADw5srikQsDEx4EvDzgmUTBAD2v4fJLvmCvL
AH6Y1s8m/kVyffIoaePiGpy6tYJiwVOaytxHAxq8zZOISvt2bhjZkPxYao95Arzy
cN1PlSVcON2AeLU5vb7YNoglfuYOJOEGirFmj/coqE1PvM2dpXEnlytshivqbtQP
eZ9Z8oObYw5nBS41JHg6xI9QWR/SdfA/UcbAyCgp+Vnw+buwLu6+KHhfie8DXNGv
2nQgIqz746y14Qh11KudTiKTpqjo9lY2obb8aDrzbfa0d4nPqj52rVqKZOX/v+yl
8wgnpUVcfCNDuH8qnc5+DZ2yjvJB7UpJOhD2x6fEamLCoTEK0Ehmj5HuRQtOLGJ2
mWohrAOkxyzvTMKyR1EMaLbS4A6QKY0Kn9VY/ej7qADGrnQBa1M96BYGKDRaGDxm
kCEmmTPvLSucM4rHeT2bP5SXUq17kg+KKPlNYFL7BezOhwKgZ7GXi8FVMtahXIF2
WUhy7ivKkSmqwWv9rK2dkpXGR+kvmWx/g6DbhraU1ABgA8Pze8K+ZhybNFE1cw43
ulDvuobn5/FyxPyMIJck3oWbLU6i6mDRJxkFIhK/wHouy/36FCEGAXWdIQ0gEGGe
gN3uHBruq4NWODcc+GWukieMoGqHC7L+I9tRZxmegfH0ilae6t3psoGg7xGdWLEE
kFeAK9D7M0Fj+MN+Scrpi9YcrNfmul6z6EOA9v5eDcdaes1wYHWWDeR3AOrKSmoG
fnnLyyWK+WTzhnROd5duaQIUMMt3tK3ZVi+5hZtnMgfRRMaw6p+cXGVm2a0RDlyj
CMxwpuYxWYNsm2cZpZ0UGQociy3iYPytci8Tjln0wbcHnSgOCjSYpfeXatWXfKAa
ETQUvj8sU532rfH753zbFCgxY5sx4Tf+S/EM6a7e7J+3oTPohvg1qN9k7j+O1PrF
XxELPxa6gtFh45yuGIhfjBoSQxrYlU4Rrk3KLotLMOjKTu/jXiFxaA68yhEy3BVS
Iszpom7R+1dWrDP/mt50nDNvuliFGQ31fvcyO+hLYfF6Sm6eFBrk1ov8esp9Scya
M0U9BkAYjVbVs5+QF/ybaFy/5XyUbolRKRtgaC+o4zhs2u4C3v2NxDRWHh1GoEc7
VIY6Qs/xmzFqReRgHnkQFCEi8kWN9bt0ff2QI0i3Fjuslfkp7j/9h/HfDQYLyyaF
novVbfveDr9p45zPdPUb4MSNB0xW4DovslzA7Qk+Crwa+hTS9UsKdqpnkMWtil6K
NWJfEajxqQRlxcW9ktVkNsN0hM9v67QL8uPFX6ZW3Zkh8ZG4rXibOoW4ReVHDZP0
AWuyKi3fJaGlphIcrH0xW2EXn9vBwZXLyx8Ct1tTsXwf8dfnIzTZYKsQcIv69uAn
L8dvwEqYxhZWDOV/C2IVJZ2wo5RU1xk1NOZFbhHb8CX7mj/QUeKMubcLmzPxpM7r
/9wcKLB7KG4gzhkBCgMG+dI7KgBIGDOSH9oLQ3ImCTipkNrQS0tcZs3vuHglyFEL
X5Hm/WonIneLSz80QaPNQnDa3gOpA4I3Cee3VZHvMJiWWd+SwUPLTyGPofxdk1dQ
f90ZyqEP0wjlEXGr2W3jWfcywX6+N1KngWTkjLoMlzKz10sVu3VoBJ833HkTwjDM
qLpuC+cQq6oig6RtwA8CcRegMM1CvSVqBw5U6XTrbEjW1S+ligW0eVApmne6Pk8I
/+nD6gK2CG71eswOwkTetAHiDsaVa5YcFMgplvvQ8pBiPw+WyahW+L0CpHB6fuXD
D62qpcsc8DL0YdPHGohlfd4e5SiS2c50jkWIjZKNDEPAkMDew6cPswF1qLMHrzdS
CWjmuA5pjrtvI06gfSTYUghM9LuYn3BL4p5XMMIELztQpcoXgSs6s4ZOiHaVGQdj
VS19LXHs2noXPTHNBh7Dch1nvbIV2ohfJjwE3q6u9XMCnsyof9gti9Uo001F81n9
n5R+6RWFx3Poly7D0Anjdpbqyiy4giJmYyw3EYuCcn3R6sW/gNsDEd1wzygW/moR
asJMfZoi8OAq5JZ3P5BhwJXv9rSCpJJ43xiHDh0HS2lx0QXnCTB9hutGNdEoZLV9
Qw10Dz8B4T3c7wtqHUJIg1xevYY6WPsOVqH7X5shQm8eOZw/Y+Vk/r3lgL9c1+mq
MgWlYbRGrsIzA4RhZ2JI/w6/kjid2XN8QyuPxwe59YtcwjXg8dKxmpFySKj0cygz
o2UGmwa184U3dcqo+XdhNGNwFLmjiNgf84hCiiXfODyb6Py5N5A06CScV6+owFt4
eWJ9dFsia5PfRBUYdfrdbpKfwU0yzndgNJ+4Zjsjr0DUd392PULby2hTN+uysD0u
Go1HQL5aPIftrHEjxyQA2hkULk8ySubUxUugcsf1VHXGMy4Ty+WWsAEuue8xqA2B
kuRBHhnrjAdzvoBw6BM6uT1/mCuRdeVxfIfbD/RA1qs47W9CjYZlwqMTSi6LmiS5
1pAMwYVLaackd1ouHpVHa1mhLt805MaBZOuuzhJT8Nydcu8stvY+Cx0kJb/3wqTc
Nmhtq0dpfTplSZSUP30LWqlSWmi2dMQ4XKKQoJ3I1KdEDPzdhtV7XaTTWUk4cdAI
VIUo1GSlF/Sksr+EOIp4x3VsXlScIgeOCIZYSbSM9Omff6tdau3rNz9L9JGAZouv
ISVaYhWsYyXPeGxa0I1smqwVdg3KVjCz9LIJSqtVto1Uyk5MDIOfRqLGFE9Rv48R
1EbVPeW6mMxV7cYnEZzjsjRbnogKbe9+hEc7KTcLkYBuvAdOXkgnDlrPJhSQA/V5
FuW0in8ow4OTB4WB6jMf1jkZ+zapnzP3DZ0dxYX38eFkLB2zyaG7eHVE+bzA04tt
jO49FujcFNBL0+uKtbaZ2ftTxjnjz6aEQx0Xj163eSNToWyeuxCV9I5bkjZGLs1B
KGOt71lPI4+VBjQW4byh3hrbYqA+YxbjonBl8f29ICo3YLXv64fC7K9cXKUVTEEi
pq8GYwAAXievAKph6vXfuyp/n1V6orZJlzyD3QsFAChGVOKeQIUl3D/+r91XSN9M
EC4XqJtxyKqjJSiP+w3gwlq/H147UMrXoZZC9DXWKbQIUiDAF6k8rsWGsepOYJn1
+zmpGm32BYOCAkc4F0cCRegQj9lF99u/KUuMnNB3FSicudn2gP/LeH1dJciliixj
bWwmmP6VS4E9rdYXPoFYR6Uymowbs2oaPe757lA5uLnzDSqxru9d9DLBBSGv+Ycs
kNFLjxMkXw+XfqEMX7Yd3Qcivq/BvvIzPOvEMJ6Qfytsoqu16NU1CO/WtfnIhD4r
oNQNQdBcJCvXTSYf6kGSyMf+asT22diDkIPodqQ+kYCn88wPDNz3V1YG2SDfJL0t
ms1pub4iIuUeA1JbyN71L2im53VwK3kWukHSJ1EMB6JXtPRVu0v9bkEVXj6zp533
yQCiUenEhYooEogLf1MROoR6AVJ8T/E9qL9HwYG24ig5mbS+fo3H4uKwP5Vqj5Eg
4A53QlAdCRL9kXlkBvTe3JC/8dCuXYGeqUeD3Azos5r2DIeEAf1EnLCgeownXlf2
cn3x3ELjJq7K0D16cGqxq6EYraT0hkHwIBRKRnIgcIR34M+blMWmgLsXMIuw9rua
HxRC5rthDPBEL6wPNDFOeyjNulfw3xFxyts0JJQRTXNqayIzmRzzG3j9HnavI8sL
uzTJy9C6sFBUqI9ORpqGiHOwBIdzYA+mnC7ETzBQif9AOqdCibrVAusE1p97G4A9
Vz2V/MCRDUe4p+NNLY6+yeQEQSdZpcpMUc/YjPA6jd0g/miTs1w2YIYgnED15h3h
r+8twcgoxtsqZfEPJxV51lWXWeCUQ3Irdvqbx9ZiRu4hkjmQRlk2+MbP9Ecl2Dac
7xftib4lYkX9D3DoFJBzhOPoe9kVBjf8NCk/0lXSadMaueoLlirwNjpFJ18cxB2O
9ChZn9E7YxqEWiC+c5W/EX/YhgRqItKeROrchjSEH+b8ztnYogQr8KxLZhIjIjbF
5dnDUIKaljo6aagXV2gFTCoy12IIomxZzD+QE1VIT8QNHRUOYeeEnJGlQIo6R8zy
Nv20dUqF7ws0YQVpyEYFjQenlIBcrvDnhuz73a73QBkqEhdO4g4xVfpu4Tr736Qj
zoR9Fag/wJCjb2FVnzBdhlGsv2JCJQWqkdPUVWVBwv7J84kr9AS8jB3xtLFgvNkM
ETOXBYG+Tq+rV6OumM6jzTNvqTIhj8baR6GUItbm8XlC8LJkXx7JuyhlcR/yMfrj
0YDuWiOcx3LDBs8xvaQ0Hbrc65RmwTQNrq69XzRTRLXDIZLU+a9YYI1OjhEkYhHP
AfkQbz/r46oTzAgLDekkzSnCPtB8+Su/EOoPeI7RlktZKdHtnHXCdeXLPPfqMB7E
3ojLUCPO11cYFruVmIFiEAdMWMKxkhW/VBKWB5BiMHtZy9VfvsOcppuSmR8DnJBp
U2oZtr7AFYJXbZEqUR1w3PeMuuDSGzMtiWSSR+38kdjQesMdAakwlwE2ilgrA1i+
k2ONZZuMjcNqQD+Yv2qyMxybgJC6EVm2zAgaiAUYJBVzMyH/r/PjPRFKzxUJt10h
ViKOmga/nzTWp2ayLVlEFJHcn+4hZKeJtQ0GjxESP0YkamEgxB0qL/hTKekSZlJU
otA9yfMQ1Jn6mqzqLXpT296sAuFbw68BHkfRI/FxORpsHC/l5PUrZloXnWR3+5ed
Tf7V7Jigx/OeunrBTZbfHI8Ed3ywo7sDElb4I41GF1x/4+95gjrr5cnTmOruUg3U
RsPzLGTgu5/h6HgQkiW1T7dc8PYymPMIXFMsonRVGKj2FLDTyTetpSyOLDWEfYB9
I/KEH+u7HNJpMhmH01da9FJTC1Y6NoywYAEXih7zKdEHfIgWnVmKenYLJ4hdhphm
328OGnsQPb1CEPILBFEIc3N+i/3Y3NbhiLEfa8BMbPE9CcA1ZNtT3LN/Cm54hDkf
ORK3vE8S2XWjygiv/nnLU6SPJ+6d6XF4pRqaxPgrCRoH1uDWgK2KHMFHZxnin/Ig
QQIPlzNgvuSSuLA7exNWzFdydzwmWZbnW5lx+/OYTfML2gVa2uWkSrceQOD8d3im
hkPA+y7XphURtbbotxNzmHfGjDlv+JArikhOIqL9BgjLLcRyec79+cVj8XAth4hI
hmf9ONH5cb+agAGHFb7ups/MK65G8Xtwy82BUReXzCGDXv3uyVqXhk5EO4Er0wqY
oNrPvqAi69tiEGx1N0F69j7ws2rnHY/pmle0sTyQG35o1wxbQXaehrH4GWNws0w0
UEI1frj1mLFmoOb0zIswEDV8sgGLFdld+9jWQU2DYbMGYSZNUXvxvCxeEYMJV/7E
4li2O24QKzohWEvaEmeMH4nNP6A/sdZuHXbAXxMXGhZf6QIJVW/D9PHkEu5bqHon
hnPBnYbnC1oM1vzKXwhpN8o7mwB+obHR/o6MeHERjbeGmFgVY6uQLt2/yWitpymD
8cjBdlNtwcLEGMpE4wE+REe77ex59Rd33eLTI+k4b2Iohe8fwX8m3e9repCxCdXP
YniG/u9KvNtwt8LX+JCVZWHafgms1zNWLY8RAfbMJB1qXl2c/lq3/9feCCfPdqRm
pUhhou2yNozvA9TnBB9HZya8licW8CAp9RWYD/N9z0iAQSwORvQbAj/9IuObkCq/
CjH4mPEfFoqzDZddMX6T6X7JPRE35gxGaa0wt6ddN97lF7cnmCH/fiir7s+zjRr/
3lOr707woA7miqMJyEkWV0eecq9qnF0AMKnfrm9RfLmTUNhIo2bqv+Ad5ngDYmAm
+AdvCVM92h8LTnn5pOmUH9/EMxDN8kJ9RMFbgTEyxp8jBIRKWb1dwjMnqjhfrD4h
TluDdBfyWBotrFPFvDkOMX5lMncY0YAWcCa0u5aJL/ziEmIoKZkcDlJPUzW9DI5+
HZ9rp9yM5oP8K3a4UNJOgjlsrq6NpuR9POXrd9KYRrAIJuOW9cmTO7AJoQHaM5UD
TRx+Bo8IdNkhxn4DYqPQp2mcYMiAGJU4LHjz6nIs3lUY1DVIQbNjNDz5RbGgT86/
ZdeS38Y1kxn1CjomDB97RxTJy7XZweYREKxxJb6TFSlE7cVF9AJFrBsxOoTfxJ/h
oekxHfpwOqRO/Jnut3OgU80rNvPTifxbw9ImjXr/sPRLymbtdBelqwJAzpUppjqj
MP3W9AgJmz2jDNpkfcpOkldv8Lcb158U7I9ACJceFwMJaFjP8XhyYAAb6XqaG5KN
rypaXoO/fnuY99Yy0vKmfXnkUYp6L6xUTei12/offl5qV+TcqsKUNTM/0kIKLiL7
uE9b7XVBiHrr8grvthkd14+p8fDUmrwixtrYVj4VlhQ2Y/kYBOUTPzrRCwourKOs
CoPbjMdGeRwNcxQ0Hf7X+eWBUIi6HWJc9Ba1D1jUoh6C9+VREMUUhqaLCI0Ogk36
jZkPyccRJWA1Ih0T96K0+QCpznDohLH0zWG12135T/9jrIWFJpjY+PliEzj+877D
Ckbp3HwMs3Lsji6fDZijopMxpKX1GYNpdAK51x/YlLkZttPd4+snmAWU82AqXo0X
ggl+8fsQYtLGMouihZByqJIC4RyL5BdSyg49Tgq/qDdwcreE2aQJkYbBljRG14Cm
i7z/MFtKtKnF93nXTT2Up2hvMJPMYQo5eaI5h0OGrssZBEemwjYEMbDrSV+DJC6g
bxVh9gyK7n/3rUMvLlKyxKSSCtgCCK2itP7BFMdTF14OPe5bUsnBpczTDCVF1SD2
GpTkG2xC63qji3vickLNosCLUabr6GG9u9H/r7LROKjoiI85D0ckw84JWhH5aJEr
pPUoTEzP4LAaTerCWJQ0zykl65DSY/hjq3MC9if9JnxOYDCbXNRCx8MMI9jm1cgS
0IQA6Y5qz0IYeS0a5bczq2+UljOphtU9Deq0Pe++N5OcLuTsA39mgiL3DNHmJzG3
G1LZbCyxiU+LR1xZbXHXzP45T5ZsmvwQBDjPOhK8RMdorGTVZ0xy9Ux91sTTCp6N
h/h0NOTjxmFP/bs2+orNIYZijfGk6uR6beVy18FWFfKAR6hgbvAhhte8I8fNboyh
XmHQGNUlbo38S5NteTR/v4utQqBLf/Dzkc881AfzB22SgYg64M/hENijtkqJUUgo
EmcNcL+uz23Mh2yi0MSG36wdT3VKgSxDjb4BGeU1MnR/JQH358tqVivGSI659h3Q
4aY61hpZ888ida9Si+vDRBL5nDIXdo/w6bYg3sazo5Y2pYjvV+ywziaB7taGdOoj
3loI66fkT+t9G8+CWqGQhGZJCIGP5nrOFWPcHQaZvYwJnLwvxgaQTB+nAO2qKzn1
sdkBxwe7q1Y7Tu02iVfIZfDfw0GJa7GiihKTJNYcMwvQJS3BljExfllEkbfrwU8R
1itX7Jqaz+UobQsUobAHG41HDWq8wgetX0FQMgANOTod5oAv8iuQbudADjvRiokT
OaV021Cl/HEqCmUc276AXUy2dcKvocy3+zIvBVAuf1TJT/raSZa4ExGz8Eq3OOG+
tKrWQGYiKG6lBA9lEAbwWpjzCLP+aDr8rg2Oq9LUsHEQt1L+ZXw2kPW0+yZPAqIR
70TVK8HHS0uDq6ZJL2UJ2iaStJR0D7wzPMzjc9Ne1jOlFfS/9kaRWxAMjF8tLAPA
hsYSPLGiK9Qnl53ZE4z1mwxliGmGn2cZ0WU4Gxdt8ok5mXWA+nyaVcYys65S/Os6
TmJ4S0+GG9HV0NxlkeQZSHtF/6csdPnwJA+mKnhO8AtAdVkgm4L/wB1dNAB0Dm9b
694EVup974cogAGTZsdFGLfNLIA3LAxIoxeFzqlRyY++c38iLOyodHXvqKB8m+X4
z8uvo1Lu7jd7PkXp4AO/TWk0xMgZ5dH1bn4WhLvp8Q9/n3NXvC6YoTz0W0zzNXnz
mCaMCAsjAQYMApLBxjHj1IJwnQWL2A/eG4UoMC3CNjxxXG1wvPnaV5+kkpUxXW4l
hiuoBD7cuakKM3MfkrKg35J86HCUF49Z6LFhLjksMaAdmxWYw0BlEypzLaP3/8rP
Mb/Yv3wcGQJQLSgRrG1SfqsY8dRncc0DXxLfGPt2zU/TZByvgQE3CNWf7QvQS6ir
xr7WZTZzrziMixn3XGY3fZLfIsWWwBX6aFe4zU1//ytxmkmfrSekb/PY6NVN+vNq
BGIvfhbYLHcO5lJ8oym8o+HfSDwtc7+dIYnJV10MRLQgFizrkls1kDuM0NgkfQ0v
pIy/zdu/lNe2UDe8DEgObDwyXP2ZlLKYlzqoKrX95XVRdLuNxMBLD4wJ4jYZqv55
ilH2OTbRRZJOevHcl+q/KoBx4EK6nINaqAZkXx01zYbWHjrlYDZT9kKpmLfQjMuE
sYBPj+V5DW498Ail5dPybSRk0EjaBF/wsu8FRdlak69gF9DsraZuEtlAbJVz6WA/
rURmTGPSgFvdZHzmR1jcWfglPc4xM9jDbtWmQ5G500IF5LUKlvn8PqDc+3ovMmNa
MygoRpPUbj3mypliQNUMJvfYi1GX0tWwAZlMnj8M87+s0eTPTXIBRrEQHKd7vBqo
t4rghJyYoK938KJb6ATiU1WoYgK+feFr4G/wIHHMdtN2uHsbHIE3F+7Wm8TvnN+C
KcYZoGnchFTLN3SfXa/Ny/xXRrWr78nd6+9N7rdRphxuhtL0vbhBZz36BAzX+9qS
nRHm4xPvD0s70lyp5h7sjN2wefY/KZpCYTh0CPFuqXoyn2wOSLFXIDCxAhEdZJWb
Hln2uuZc6ZdPAdd26DnMH/rmlrgjTWt+rKjmvt304mnAX32bClFpDmfYrO1YG6Jq
UP/agHEP3g11Aw/L/UAB0MUWTy/JcRyT7Yu3FuMlKYvFmPGUODfnoNChC3Jxzfom
ItfahLSg4PNCrJr4Tip/OPZV1UgUwFmrlVttJiY66QwxuaCFMEJOld45x9hKbQju
Uax0AMPB3qRPSaTxSCRvvH6+cXgBuzoapBI0aIz2RatJi2sxQ3FQVlsrxooTWO4z
voSPGLUqDdayQ96nPP9OfOHPcJOQwFqZ8FAWnI3Yjik8E9lueLwdTQjK3Ti9m/ue
sfu0u55MhDfqR0CBIljwjeRFYaDPWZP55QSNh5nXtf6DJXwePvEZj6oJvwTO8Ts+
GuM3E5e1HH0HxQzLpjXKmTPNNulQ4i7ZSZK3hhGwCWHuVFl409ymobb8cTCF0MJQ
uC91lVsD+biWLEGGAq2OD6U208tkEBZp9EuGDkgkT+URrNzWvWAGgN3ocZyOT6Xb
gO7Ult4/Csx/vKjtCkIjCgb1e0iSEdE3euG6bHQ/CQWdmCmWPKQxNup8EwsQbepQ
vLuWScepp7/tB8X0tuHUXVcXCuYBrBPFdPJoFwhSA9lbBqQjw25TKVk9rMK/c3UG
ubcEEeUpafnIJvwkoFTiXruositbSNz7axyDnTPWJQY6U0ebLDNUn0pzbohm8Ff5
/hoENON4KNXCvEnwVq0zW6TwU6IGLY9MX54X1BMeSYK4/bheZM97pCFfXjk0Fsr+
vfUC0jjBy6uikE0XsDBfpF1LYcaC3KrrOrUXjLWIG/EGFNSkK6r/+u5cd8LKMg47
PG9HaT9sQK0daqLdzaLrs219dKUfCJ84aBNkHPR7iJSL/TDSh0w3gMRlmX/FOY75
obzYGPo8/w/RUAS0a7mOOrpNj3v1tC+ohp8XDNtctljyvwxlwyjYJlUmEFMvj56W
D5bNpE4Exoay38yNH5uhrYqLJ1jHAb97gSeqQPNiupZ2/D5wGPntGO84seEgtml1
AnrP6EjC+TYfyQL+EZqKImqcsbAkwK01uJdGwJCvlD4VefLJ6xaIKcfyWo06skr6
BO9I2HXPzNWJhpSg2V2oZLkog5B6cUkxZ7V6Xa4aKUuXfSB3YfX13Y9iGADYPL29
6pn8ttMh7EdswxjQvrrw0m2wMvNjqZ8JlWjDX+siDV3QqpOlirQMfjjS9GlX4nlC
XN7+OvPsFGMLnXYAHVcG+GFOsC5IMCXIFGOw8kKkMxl65Hgnn6rhJCRy8+jR+L+6
uUxHvKmB4SsNZ0MU0w2cmYB0aXI6A3JYGxb/w+ank/GSljVhqucN9mr4BVDoaXEZ
LXeuwpJyfyKt94DtbZB8dM4O07orqtW65G9B3w3MkurSPBphykeVLmy8EUsq7txQ
4NUps0JkNWI/We7oUJgza4YwjInIygYvl6BRZSDZLnMEy2PW4nw/qYf1GaqEFOxk
dKYg+EgMhC1ZEDjQtrGkGUKKDKxf8DuknotbPJFE8duRViBOq6Gs5EX1q9fuoVes
M6PVGw2KBBIosCx7T9e/4eJeQGroY9pH70U6ol8yI1v0rbuo08yiDcIQSOMPLbnn
hiAt21i4xFcAj896TZYbUwiquYj7fAEVczI1xlSHcm+ptnSSzrzoS847aBtvmeVy
iaSUtCIyNjJToAGolwncCeiTNM3z0FXrlVElSTbzAa8J0JP8lslnsQyx/v0ljPok
kVI+9XrlOh9sigWmd2BXL2k0ouW79PwiRjgYxEGKyN5M2VPbzAahtPPwMHK8vAWA
qqYeMn/R/d0hz+E7h95YvLzIX738owTRkpWBK8ExqzHyBRY2jG99C6GI4XuCbx1/
m7RhKerfLYzngynnN1AAyGYr8ZLoo7y2PnbIXYJ1XZByv/847huEOFd4I0P1HNsb
cTHg2Ifm/+W9guCtgMCL1gkowZrwWMWqDuFyHwb4Nmj8UUWkc0pR9bCuJoTPlv8b
4G9j6E+pxKt5mwEtbPWQ+8glYD5yzkA2K4xLpy3Saj59PZgpA8vn9AoIPKrTwLV1
fmfuorfHjs/peZ81Uqr5YgMdASINmpvAxa6gbNoHgJEbXXyso3iMTe6Bb8GuqHfF
FAYPc0TCe4CbkGI+oFkIVj1BaLcxzdxXEkVbB1gkthZiVVra8j3M8NgpZVd/RkKb
bV6jtFdg/sDTDgHiSDnYpGDwEPhc4Pb6OxmMVDSrQCCFhMEekmQnr2Khpe/da/kX
ZiIET5aIK12Xs9F/C1asw4u+urCGCCeKXYa6By7srJ9DkWpzf+GGRKAkUoWmQzZ3
XgKaZCplFNTb202jY6VYA0J+JE1vvevw2g5p7DUy4hfzn66pzX9FsH5t328n1Eom
TQ/mzvTHP2J7En6KeggW+Wi+55LoMNHsTwsdCrO/jC6pp7bT32ID48V3l6gqPx4j
n7BeY1r2l2fc7iV57rfYWnekLcO2TA73EwW1/zUL54UGcrAedW/wSwDN2EJZLlK4
tvBvVdPKBbE5UbqqEOAZW/zcdzMyHMmScbntQAFzx38/rQ6sqREPJhWOFeKhRXQf
ur5s4S4tt3HQf8M8xsCPYmejgzQUvEBXoHHZZQ/Uag5izkhXs4le3eqcgzf+BoJV
`pragma protect end_protected
