// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:42 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bx5jW+mG0SQNlyHn+F9hCtpsOEH20fEUWkPmDSIpd5tTeDLqilz19wP3B0xRxIki
bWPs/A7Jl3DeLXbkgPKz+CT0OnZlTc3lk64+nGj1aTMzYjTbLjanSfOMT+qX6Qkq
jr7zq3jUAICe8pEOxCvV2HxUtuthNUlHlRDW1JP25YU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7104)
FURy74UdWyvb5xVATF/fQMpwdRc3DPGA7mNtLpnZPQH+9eGaDiCDIrRTChzrlubJ
0+axEOPSklNAifyX56PIwB8ADE7Cne4Dmucgc8mF8djD9J/yvYaEXM5obh6J5vWu
yVPrb+1AnkHcpNMW0DasE7L6eLdBKJOFJ8EJBXuD3NU25+x8MaauX2RDrFAB+0b1
yBhQ2WpOa2hdXPg+p45jCD4Us8RVJde0v/k3uneiaTec/RrvzmzwkEF8sQIfPShK
9yQBQJCVhzGjOby/m00pxhGn8Skg5fa0nRV3gyiS6yB4eAhgNmY4GgDxGHXQUls2
/C7qJo9rUkovciTIimvym251zxBRn5MkyZBTnCPNnkskYtgDIyOtP6d6uXwCt3BJ
YQvASA6uoj7Pb73Sh3OKLxK7l/0h7MuQ+P74YsTcEtQFo3rDS6NfxSUDkm7tGUEo
ZlJN5uIqcqtzzKzPLqrMK7i4kOfzMCOssxg/P4iIILuvalBEd/ISdyYZgnqJhRxn
wNAT7xXRHoQ5kDoOSTXOGLGhBaBIXZmvA44KA3XgIkArsYsIDfv1qXcz4ejtSd1H
Gsp8JEy/Sl8qEXsleJ9HqDEp8r2//iB1V5XHqnhgAmLPAhFLDCSnutBEfNxQCv1k
E5SvSf3jDBnobsSn0On+vQVSk3PzuWifU7/lwxZBRhSxX9aqxndOIMiZeH1Co87B
PWRRaTnNYvfmXt6VtNHzNYBOZq8enrvDCm4R6ZmddYjbOaG7d8Gj9vUAPyXYWdPm
7uK+R1nu1i1exy4RF7YodUvvCOaGpSrxwCaaD15BLLGSs6YMD4mYIskHEiYp/Tf+
S4MOQYDugJDbsKNQXzgeEAnPEpbD6p3JYm7j7CqU2lMTTjicA3+xwYeMa9DCiwFs
2M6UG1JyD9DKKfXQMZ1zPfYPrk1FtDFMSFlvrbG+dY/EHGlKw6XbAz7KEo1l8HfO
NPVfSGD6FEW7ea3EPhQrXHjqmJon1BnKI3Zss4Q8aiazeQVYcxtzb9QZOl7rh6cc
l7XYJyG0mJHtiSgubBEaeFw2nCBx8ek6R2eNIVKm6+yhkhIclqP55whEgiXkWwU/
b0/Kk8La+Bd82ZQuehI4kqFis/bxNuF9q2t5IhPFXo6oJHogGyo+5CaW4VT/Qhed
TI1oqvhumvkz6I4QLBOB1aFShggDcMAkxlFqD1d6ozo+yuYZcz9ExYeG15QioRyH
ENezViGqp8BiEBIBpTV3uUrbUXdFqjeu7r3m/2YgpqUd9M2ENfrdeYunfyGmHC2g
8q0jOwCEE4dUXAfcwYIgL4jUOwV5v43FsEVmc2qCnh90zV69pEMDevovXcs3CQK0
DEhyDWuupi7BMCe9TCbjczCFI5vIEEl9Xa9RYKAZzVqLRrzK5T0FcHcCLLXY00FE
rA5MIqqWCOXQzYZeB8fHyRf0thKVRPbfuYdJwl+hB92G0U5Ha+pzc5e2peF+zaZL
UTnea0ns1ZZpx6FOlkH0vlxz34jo6n6wT1u0NK+eXu316k0Wh3iBoQCxdaMY/osT
kUHzQZFJP0kpnxrIvysmUgLC+bGjaJOWg9aFmJ7RL8qjsT3EcxwZmAXkqK+ib7JN
mxMPPoP+cPKdAG9Xl2FX+wZEtSOVJbc7ZD2EL8s6/bO+sP9kgSuXYcIWQFXjFkwK
sBfBOT40tefhXnVi+IOWhpdjksjMvR5W2/9lTqrI1YDAGtoA9T2APredicpqL6LS
3wFTkeq8XyAwUgoR15f8G9vN8iKbuSwdHB8ADSP1UV8iFstvIrwpcCNVcc66MoW0
qmXt0M+46u4fK1OvSX0xEhG0rag0ZZxfRBhFsXvw0LcYqFCuBpJcuWFP/UWsSkus
LvMWAamXs28BHxiM7iYOLPl7IdrvWA3dTy9295wQMVjt1OOZ3lNEGVOE15RArbZk
Cc7jESiLwHbx0AoJYH+Zn/3J8thz2MvGmq0Ob2RoYA0D9F/vX7zmZRyzf4tTSO1L
dvtLvbkmbin6U7Nf4r290Zzj+IB7bLbjnIkBCiV56exo1dRpZuwb7PVM7xxly254
zjWgSHLxTDzWuyWwpWHZF1zRVTWCQFnMJa44doqBEqKDivpLyJ5M/U14P4c9bgJC
8y4ucQsvIDkM2qVQ5Aep9AOxv77YTbIXMofEr5HuQ75D2nDmiH6MXvs707CDSC3s
KeEp3/NbSTwEpmLpZDtwLlPdjXUOD5czRE4uPk3UnKfyOxtMU3eHw4hwAi1HVAPg
104GU2bchnXcHOp6/PD+abKwsTrk8eGkHxtaqPYNzYx97cU2zNDKG7aORlI5MkUm
uQG5NwrvmUFtFUeMD4Mwup/CuebD4wIXxiS5TuA8tybJwoYt8CAMwE91F0t3INB2
PoAIPV3e67s/DVtiAFHz4KZwWSiCA2guzqU8F9bCwvjcQD5o5O3pv+ahXA4ONgkA
wpARhScYbu70NxapYyGvgUUWYAFVPo1aeXJ0x3H6poFdU93T9/7DwIg6jmDWpLJd
WghGgDKubp/OuWKHYWu93aOvEEzXiXjOWk0gPaiRgQpnZG6Qy+gwIf0eb7jHyl7J
pi3fEMJrQa1IOVWrqUqE/3gEulRBckDnKUjFuDCmOY3daQxI9eQvKVyWpbvIRk2O
VUzkr4F3SfrUk1hTVJ4JPmQQSyk4hN/m4QEy5naXQ3VEDbv66lQZvdyrA5uWhu4q
TgH+spDj0z4+9dz7oIdhw9go3ygpzHVWUA+6h/KT7ePSG8dETmoasyjR6krnZ55f
+kMBLetlWlFzjxDGD8cocOwDa0ZKokMusrLJHAskmJ619ITG9tUgH3RtOLXInEoY
zUbSvUPwiUXeJ2tZ9FQ25gKeBSUkT4DHvWNaKx94JcMUS1Db1Q8NZE7e7BcVWIMj
oMippsEfwXMzwygz4gfXdSNjc75v+YSoADqflPsXPlqDuqeMl0+8errR3/ldkTEy
r3KP3AFluq+ngsBOW/b/d5ff6q9oTc60KFyoscbib30K/zegAYPd7BmTD/+gxIIy
zU/+iaS/EtMSmhHQdmtjzA4vlr+2GHRX8QyawBLTjjhalcb77b2TKPptUJ1cxOGw
0Y34n8wsSSrctNSUB7RE2KiW5MGWmK8m/53TR5Tz1PynQDc5AX5gruPACZ+pRZyC
2H3934Eco2B1PGzriIbA3jQdMv846Mw0HUqAiLDNwWy4oidWnUa/gQQm6CNeXW9J
2E1alkAczJpfJMVoN8Hd7LLOHWEubm4YqxVT6Wb6h8K3aC1t/RwQ4DUtvPGGregH
aHe8qj5xf8m7JFvXn5cTGLyliC8DLyvjCG/CbVmWyPWpUwY3qiCP9q5kF/n6Z7m/
frEqmGB5Sab/d3ifiYurRcR0XBDs0JJEqaZlTVU3EilnPTpzg/7W3vUxQimS7J8y
8GnSk5buf4/g2GLwE8o9ii1ZrWg8C4db2D/oYLepYH31/ERjeR4A6TfWpD8Qm3+B
O9p/+g/Dt3wdLW6YIn9sjtFigG4pU3x6uNFz/pQ2gAsQ+YlkHimdY0FwsvyexJPQ
baQfqKdvaHuHN7ktWB1OOtvXvitBq90Xkux4u83DMCr/PuEhvXrEjhBpiBGPVIC7
a1N0c60Rbk6lYEH1at4t8FBUTeWOdqt0lw2RDFk5Y9qt+4wVHqdyPAaitL3rJ3a3
X9dKa2cQE0F/Fv6hRu7tO+1NgRpyspCmdDTOvITGokVHAIpaemxDGraHEYZLaThs
w5iU6fjc//o8X5CWM+ueiG7x03Vx3ynhKiqdLbfWzhVOEg2bw6xaWYt5Qie+1Cto
4XaML+CU9DTtxpQmtO7UHejluX0OqOAvWYou6Nywh7VOFBMWCfsl/MDFEvT029W+
3WvQgt0oikOjsXR4kznR5cx7fDNPZdJoYwm9H2opkbgEOOviQjFiOmOuBYIohq28
FbPBAzHxDfWHsICYKkXhFibAe8DsXpkiQBGo9ClOpdt9phw3YM9F7zamC5Vxc9FA
kODSD3yEY1Bd6Pt4nBxiIgxbuNq2DAajpddYdPxxJHfDVP5cQomM8lHIJznMrj/8
SCAh6TdNDJYTdCVJNt3pxxWjcc+p62Tou79ucxBFHGBUrGobpnXLSYM2HOTgdZ9V
cadRQT/J5y1tAtrvGjVsxTACZ1Vxnmtg/+YdJ7b9913G3ZspZMRxGE8xvWR5NK6B
0f+PR49HrWAqgLhw2W/ym6Gjf/Vyk//YkctXnISBgPlqCIwTBdt8tUIYkUFQ8Lrm
2xbGQ2t4q+XeGiJJglUHEbqqjKcW5gQasyZszKE01TMBiAhWLK9zPqdi+ZgCk/4C
PwmB69UbotzB06mYXDS4mgjdqwavCXKikQC5RFPrhFLPdTLZ23aApwAGHletROAR
11VILSwJsyFQzLXHYpdv6cOdkEcp6qu7df5XamoGJWlRVhvMYJN5+kR0WlIocsh6
gE5zDWMQU95gQvec4QcD+0w4HWh6uSb1ocZKYidb7BjIcEwB5/mnBFzPLjU9/QJ0
uPD3vaAEElQaXKlBAXOYk3S6wz/C36SuCwrRrsYO2ee6zpBlize0IWfIK5XfvBIL
3TIVpiV0uHGGCjrOXAd4i2DfFAQvwZJATFJL+aMwYw91QLqC/WIhAicV/aD6giaG
e3JC//zNHS0r+hEpZdubjJhQjqQ0v691/UT+cMuhOs+Ki+JweIJ3yIX5Wy0Vhtei
stM0ovMXXCz7Q7QNZ1lau9gs/WTERIIzAvG/Cg7ZUIk6IlGNS2a9//QkIEQbC3jF
Lp4xfJ+rRJBEoA8CXMqyeTHROVOc06DTgRfQX/4ZEsItv9NbBHFIW78B/+rToUO5
XHQK30h9eZ6mwSSFmKCSu8fDJCxLxe7Ngjfq0+SzgCHxs6dN29VaE1fFh6T2OhW0
piAN5JoiAIhmFRcR0BW01m1XgCwUtZrXk6o/29cvWfE6iZPPKnd2F09yAxrZhS3v
9bYCfuixcr73ke38qx57iWyOBurjr9FzelIwkrXs+0oEa04/AGZYWHTnXdpJ6UR2
NCZN58zDyTgydbiB+8ecZVYDftd+StkWy4u4QZTjdYEyvSMP9NLbWApfiHvFVUPh
c1LgUNWmTmP0uUWmrLAcnSEiB9Il+KCzhJhZLs353gGwzsoH/qzJEG/IdS9e/a/2
ouYqBej/O8lqF4CoGkDKwq8z3GRJiT8A1Zvf6ODetbM84uFCsDirPm1sTHf/Wrbj
y9oD5fmRVke6tvJGC++wqy8W/RAtGVU2F8DdPunB0Noe/B5U9aV/PbP+2fNH+mVz
hUzAqOaherZZma4XqADn0W8z0kMa4SmzybNWNw6Sfkjvb9Gb9KZYpyUSzvSxaRM8
C2H+ZccKPPttMuFmXsVwI2sZk1+H1nt7JOfVfz4inDtLpBLipiYyF++IY7+s/4tK
+rve5I3iBmFf54U7Ltmib4NTOozZrAEuyvoGeGbQ50S+zbIWhItbgabu7PhoXyyu
2BCVX9411y0KqaZ7SwxUmML1gdZ+lZUpTJfomJu0NPSg8W25GeUNMivzu5A15wjy
qD5GiXfM+WApKyZLen9fTq6O5yCF3Mj3XyTreD2kiJwtVGZ4aiQ+bN+1ALOoYgRg
opn3xYz2a2ZwmCYamiyDfkLstk3WYBjOrYfXUY0tSz/bo04p1qiW/K8mrB5htbVw
mAy1H4mPr+xKbbB88Kc9n0Z50kDLDsNbosYptnzirmCaUtzdh2OQoJJAvmuqttMb
UwxismfJgqW+2Sa9hBxAAZHifiK4KWnBPYyPIF8CdsKxRnvOGiiwmrzw8YLjcqvd
MEPe8YFu67IlVdwrdpRLX4mz+vQ3uHZUx5HnG58qdwmCaqzy+PgHh5OCPLayiblu
P3VLJ+kpJyPUTLDES7xZOeYBcRC+y9YY/J3BUUmv8XzFqQt0miSGS5cuOSK/mYQD
fGX1AibsUCPz6OB+LNl9pxl2bVtImMlI2+8vuSppNl6xdRwRc3If5slUhSrLT390
ma6mNGae28NUz7JtPNGG2Kh6E0wj2b1BO4ITN+kAbjw0HpIbyEYZCau+vjkGEcZm
oOo0iCU9JroIPHLws1Rxr+zx72gfFnRqKVgPPb5eGI2xrUkclExdtDqjGCRgaRNx
d9nHwjJj41gx9vo0LYwvaRXEg4b42N2bV0P/BteTPr1mWrsQSt+Mz8lBEHiixOYs
CoQAU1Dt2tRGj/eQj9JQwi0/KkN5jzTHlzhqekjc7wW/v8pJdxi3d+9+AlUMXJPm
tdItR8N3NBs0KvGBQ829o4FPtM2g72/DQFCUZ11znYX+Skm9MKXT/CmvBzasxGMu
3GrGGu7ahyj+kxHzEE0f01zDXVBHhAfZ1yxqV5sR5P8guxK0U5opf5rEcvxiECKJ
CNwfifkRyzq2EK8Ktb3fdvyKT0/RIHZq4+1C5AqcoMWWTXzXmkYZWu1uoTDOGIl5
vCo6bc+d8c5IAGqj570KMkYwt3h7xArS0tyJm43f4l3dmYT9J1haz4bGQpjXcpH8
3bu7Dtegu/K0IGk2mKTLwYvMvt5skNthZ+YVK367wh1pl/rDmG7N9qnIpx7T+cGN
aeNaY3PGLflMnnacilkhvPR9rCR5LNWCAnRgrjR7CAa7gMVzOwRM/Zl/rZGnK3am
vhBEl84CH3UORtORQjB59hfy+hFkz5dWeR0WygDTtS4tMuvgJrifthgM225xOAi8
lxjKT61rxWJBk5ZZx9W/9eqJkLVU2uOQPPWNM6WUMZRymhlOMx1GfNgmrSfvhd8A
7UfoXL0jFVi/CZCXhxUqAHVEt+azNbv3QLiuaBgoN1Dxkxtzd7urnpyhEmBPEadP
ZiOgOBHoTCOblywTUkcV68LAYt8DHUaJ8kNW8k26FKiMs8JO3a2XkLD8dahz7gr+
udsiHv//SxNN2cgPLVdUStwJtCB8a2iq4Zi0wIx6lFVPbC1KcBGb7paCJ7sw+XGj
6QAlZ+KvSvCDhnrrq3Gf3bCitPlEt4LBr/d4oMyorj1LeIjwligugYRy2+fbtFoG
FoEHaySo5eBDEKCVkVldXT/wi6HXtBNgzX3J3edle6lYORo5LymI26bgb4gj7Rd4
nQfOEkG32NC6PxdrIfEznfemIqb3TqKQaCteSjTA8lj2334cZ7Tu5IOPTOEnGUJN
+Fgw76vpETebkb4hdOuYBhColVqIGyDL/ihIO8QWQh62p6nElP0VdDK10U6vfi6J
xvJw4yYPmNgGDkHAMgwYdfOZ0PozhXkcuvjlOKlLZA/q0EOFQ4WqTOVjr/e0H4jr
SwjXsCsPYQLSjGg34eVJSTR9Vqyf/BLOZTETPKe5nme0J7YtghyVSZJIJJrG62+C
d2c8Qut2Q9uLDWDIWivZGrObLQvzv9/SobNwF0g+DEb+tzOr/ZObqKht4NcabJ2w
duJ4Hd4JDRM11IJxSM3hzLtAvRXP8NQxnWeJ9548aFY398B71A0Fe5/yYIVbsH27
A5Sx9GExswQQW+Ew0u0oXACH3sxEZAQEobw6oqXkf9Rc78fx6FVzqD36MTx523Of
JlEBIV+CIiIJYIsybhcuXWSgrH+AujYnsqeqPqzxOSB65vmv6ETyK1HZFdU+YZyk
uiWuDurpX+msZ4ZsXzOjq1OsjXn2dqNn9NF8xcciJEcRQD+J31CWYxv5br5GWI2O
RIC5I7PEbuk9jVhrSdUV++DW75uLAKrYwByXfFr2X5L8RWepMztgW6vxHvwmmRst
upV9s+1pRlFD8kBYXsghua2FIbrWUgI9UGHftIDk3JqWo/kxgd4xuZdIDvrcrFZS
vALC4QmzO70cnaE/gFuOO3Wdm1CvTH+jCzX23IedFdthfjuh23AX3TsduWkgLFko
XNDhAfW+JlJ/x2evNbM5qX7QUshjeNZRim/s57iVEW2O4vRTs8nGhwbjjROlZXI5
iCcw1RgNn1+KQdxXIA/x6eBjIsIG3ZGdSLOVHGGQ60rkmAdu9/NXC2rOWz0JK5PH
HyPIaCsUuc4QRCxygEqUhThwREg/iEKusCOBWGdmf5zs3QyQbzfNNoL0wvQhSKoZ
lDx5sHxhRryxPLhlqhA699rR3fepaKmEsrmhlxeJMxLOWok8cFutWWFZ2jxuvHqS
Ckh8Itl8EKOuIu27NszItJWJZ/7qHpkxpEwrPot6ChFHDsCXjoVTKsV94j9SO2Y1
39OljVKeBcLzvAfiuw+rrWD8RxD7xEcUOlJR5c/y7WV+QqITcSQJnAGZPzzQk+4f
ZT9MK3LrqOq21DhQn3fvmusKw12tWjneezL5DPPmAxru9EtYFAWp9i3pTusmoZ0X
tL/Zp3TeHb3DDba1WBT+1O2IXDbJy5PyoDKwo23uPEUhqMGNsspn+jWgf7GkRtQo
06P43gxg7Ku71cKnMatCR0wD85rwbmPR3i5538CZPuMl1Xp7+jpg+T1a5JGSQ5fJ
ZcyU4YlD050ntJPqdFb4J41FgfjkhKgjVEj+uYw6bfC6lkAevggpxmfYrSBpZW0m
strh5neRXYJIK3wOazV2OV3yXvQrQeveeUOzQfC872FV2+JFGsd28iADLvdpoB7+
p/5Z6OxMoGEawUL3a9UEbBwC8tkLLrWaRQZw2rxf9gv4S4iLZvgv/TlTT/V9VTuO
XxuVW6rkTBzAnQCDqSdWuheIoYESbntNf1r3PefF78nWq/3Hyga3mY/OJUcXv5ry
VhTeqyHvG+IgC2eSQueiy/V0bz2VslSsBKs1m9jd0xnSxfv6+Ok3U6KIIn0PvvnA
yEmJr/msoAPjDsC41AYYb12RWxPuVDdL8chDry53ZgPb6QDo10BluklNDWw07qsr
n5rzhcLPqqHIV8z14gD5k5hQGaVT/oV73xjf0qGrDWm1GHp/gSIXhJveobyuEwS0
54FsPL2ikMyOHQOAWfZsNzaGeexffSM99qGH5St2P+jVtoShyDMuRIN0+vpy32QO
dVXLQAnIUJH8G0njoNtenm5uznn3uFJTU20R5IkVq+JemMaX1ZKhzgQYFsvvRPD8
qk1GKXS8oSkKb8dFVxUeOzgXXovcJCbinPqJeGEnqaLMOmQKYGxu3atU9oE7+JlX
pNcDsz+BZLna/UiB4U0hhnoEQPGTpUPNLckkbdkPFQHCTLO/QwWuzwOCzg39U+dR
MC437hc38FrO4H6g8wgGn2qYk2ZTeUNsYmBMaNGOf+PjzDSj1BV7wG+GgNYz4Vms
vQ/AyninVxl+rdeS6f5s5kgFK5NrjHR4PKSGYhYws6anK6gKfZzyw3zWqq3qsG73
f+7/ZfMJLX7yrd0pHVzH4+ltGr2AdypSbUmTxjdFDx2oyKSjCuTDvxd+eKTBrPyX
vR4CQcjeJN1nWOmlvc7M3T8lUUQboAT0ZnoFo9ik0kz4/dMiJpwJufOOsAAToX5y
0cD/ZiwpaHS78hFTv2T1jy6ubpEFViPIbWQXvs14Numornv+IxfeuNsD/I7k3RHl
JAP9YN86Io0FdfHJOILXPll+VmSque6WCMUteIEcCYvC4R9adBl0XRgvxSC9ZGXK
`pragma protect end_protected
