// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:30 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ARQHDuUcI3JtDHwk7PkVjdxLRzo/Y5AwKaHn+kAzuRTDpIB1J0VTBJpCI0lwScxD
T4j7NA7JFZhwp8wEEytefu4GApaZ6HitbGymhvnIrEBeyKoG17eYeaWe7hDp9NPM
/mV9aFX1DTupvivareHox0ea+fqZRJ74JviROIoPItE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
ny0s1dlygQFeuePl1z4OH4EGz2MeZdXrGQS91RtkjwoN7tTkRu3YIVEUlabFKxu/
UtP5OX/zs/Omy0Rvv/V1VjSrEznjUTxgz4WM0UodXiLOJ0qVOhMkk9FohCyyO4mx
rAgitC8k1/uDYoHlcC13hI0RUeFimCEi3k9oBHJWnTsmXaFqKG5XfS7mKl7IJ/Tc
/Y8rXAQqFKwAvYSwURELrkFbetUMqsxGiMaOs6kT8qv4xBTac7kEO3MQ57lz+XgU
h7p4DV2Z0hmrKE5dNW+AlFUguMOD3zIVy/Z4dSxQa+Pofi2DA4YrdM78t65R7qiD
MfhTkupaKSA9LNFOXpy4l1JZlj2iy2M1ZffV7hcwhiMB+R1CoNVPqexci++0t18X
zLjO4sdvAfYo8FvUpitGaPErGJkYUyKj7YRf3jcKAOgd8UMn0NDwM8b8emq1gN/A
JZkF/SgCUkREK+5G5gKbLh7ARq6gwpj5agcZNAM71y2aiOjlkVg3TjH7lTcc2u4K
67CHxnFmlU2EEjeit3EEj58nJIdHnd1y2olpJ2lmcUiwr/Oe9Ln2RirEtJQNb0+1
y9009WhzTnCBTXf/Qr7dTRgQKwZNgg+XLoUdgK4BgTOkBhuj4Et8+qKG9w/2tlbW
B+4tMehXXYP1KKw5IliSj7CLQFBnBnWWXCBBtmuPOzv53s1uNKTCXvCeVcIHMnWj
XgJq33o4ehyxKSRYOcJeAC6EgyMLK0J7u9mkNEqY9brPHOUUtNkAD/2vh/NW+pUb
O9TUaKs/T5jBE4IWtf8BPN0JUwkK1c/NeL+Q1m98Zpp1CCgzY0Z0qZgHAPswySY2
UDhVmHAy8ha8DBb+3svrm6ztl8fjmtMSdwtYd6llI2VGTPTWHToV1BwsUpEKFcgo
olJhilTpgl/LjVs0tprdUilR6Zafp7u3K1O/BY7hBY6y1tKUNi4+rZ5PCT0gI6p2
btHOssZpTc7/KFySwOJ7Iqr4ALgprdNHyackZf9dXGVilbM83Aa3vuIpXv7qSBhP
DsTsNrVha7IWiHit6qv78CVRvsivM+w05s70p7DkEV2Knof4gA2mJd0SnC2WsxcX
8nE9gPv9vIlJY1+iNOiTOvks3ya1szULSsMT0xMt89Kc7Pbic/B0XIpo30lKXOhr
u1wma3KmRhJiye3jryd13Cid5sI+tWUuUrg25R4ovgG8Tnb52S/TudP/5s2cshX+
+7beZDKNJBLJoPIZ5C3p1XDePHI6XsL0jKHOQ1N9/cKm5WJ+mQQyAPXySiR8dET7
SA5FgfB1db3FYWwqVZ/7wY1Vy0fIn68BYLFU0fkE9TwaGDUBAJ1RyRHt5wROCf9V
5GyVye+TBFzpL8Y4VmYxaNxBAwbAySRyjGQYCKzuafWCgw8aam+1x//pfHX66Itg
whLejP2odjXMovLDzTDc0vrvzajh6EjOf3/4fCvi+w8L6uhgF4ldZPmb6ySj3UBl
rapTeqGjwT9GgkmdUBj6Fi4qJrw9q3gqU3lRlaOfyoY0H3dXFoPjX3l3kSeFwRaV
2pg8Qexcb29tSBeTVa+cVLzrOLeZJWsE8YBse7QzW99awbF/SRotjROGj24GBWq4
qwD36Wfdcv5WgLROuFlgYmUC7EwO683mjRUb+Na3m4j/BFuL9miFIoe4lQAzKm5G
Ar0rYKGI/QP7qfFEFStV3ifE31PFEO3RRxwptPURvplFVJPbS1rPAkJFdgve21Mq
P4qYKtKngdBC2rLhghZawx9/GT47oWxRfmt+Dq+XWWFnGzvJlpMpG8MnH3P9XJbh
64P4zhm4mfSN4IGzISRDUll7ubfMwIvkh1gCcbJsMsXbIgURqVfoxdHuwgiEqxht
MMHBg45QepQFh8fzxaFYJG2fXjzRwkBgO1X0ggAI5QJ47LVMw0UEtkKG6Vtd7qSX
yQVz7UJR+RorLL4iraAV9ZdFLoIMrwYjZxCDhgfrdY0pWIuW1rX6luRcCuS+FWKv
F52pdeNDYkBKHpyZ5PZvVxsgn7JRVX+ydsGHPkmiUZuA7M1zOfSGd9oakt+m44X9
/YJIZwXTuKC06FnPaf/2LQHWvMOuL6XQ65d3kAHuQK+IwPu5j3Fu7uK1ZfFoWiK+
+uzoZ5YVpruSh/viUcTCjv7p7zWImKVRXGO+ZDgRdjjD4rhHev4NFS5kvRsVfoGP
DZU1TgkuWHIx3SvT/dTJJkYuz8M6La7ZQrIkBrECC5QyNp/VINBC0r4CjqWboxCj
gRzLwt9c+fILTHnI2JoQuFH87zDc8O+gKRdIK6vjRglB6R2CIJ0ZdOGTOtvpWtxl
8jDTD5kFWrygFCzQ+6XfRO9uZvbj676HCDj6UT0AzCKY+u7Lwi+qPAJaTueJEbTQ
JA0t7uAJlmdxZWfxcTiHIqpzYkPUtJYYKdSFnGWw8npb47kJnCfEdCXhrDuOEqsl
PBVGWwwEOvjRWN/oMRrQxwzWsj1GIZ7+D+BHdzKoOWEdtSJAvl8O76zbfkc7LpVy
mR98XkqV0aX0xDz4XU0ybBkoSGn2wOQbJwTKObGgtzueQ+KLT272JLbXwVnHXLvp
cmyTwcOs9Z0JywJAwBpCcdPuDV8rJIYz9QQzF7CzEOSMyAFk1mnM8UsAsGtlOWQN
YA2H0gUWslAZVfWxqyqbAVPS+/twfU7JGj7Msqlvs0HdpTSb+p7OvEteBeG6udhf
368wZFuJ92McwkCGulEhHsuvlE4Nco/cmMCdTGYatCmcZyKmZur+RXuYuxtYTtAi
ATDTV9rSAbXK8/mgij8kjbBo1Mleg5xiHmhu0liTKi8r8Rau4x3SGxlVB7JHCofw
XoUlXmXyvf85UtGDb0yNJJeirMLqn5OP7iy2JKCgPcB9gwvszuLg18ilFsVqJSNB
7nwK6k5wM4/AWTjrjb7BqvFZgxyyMgP8B18vjmlAzCk6hFn19mQBxpLsD7NYHWmt
i6+3NNkk1NWShQWhtm1NBkCsuRHRwYzYqaSDKWfIJRyw74Rw/mzFl3rl0PUxNLa4
0TmLypHMWoQF9H1H9cFury0XDOG3b7pyEANGHhTqGAyPrz4nVUMXceLD33FbAdOO
h0qF3DF35Mmf87nNmx8Cz7foFAPkBNKTwlB8Zo2E7vk8VpsRVvFO+ORxBBlv8azq
JfE80RDb4mSc4sKVMo2PtEkK1Ub+4IJHlsxX6eULxB5YGl7eqS+kmZsLN4GzUY3u
0tT0n7RONXXvqrn+xyE6LPtaUFi0MxVALSsyqS7SExJQWHFUaGcS3izOdlT4Y0jf
PV9ptxPbY1LJ5zrHLubDnvSNJt4aI/Ywl3c9/SUp6Rtd7EngTP9BFHv3ArfpPb5o
ZHbSWW/0SxX3g4XlsGnQIavwe3mcfP08JOvAr+DRyawFvmBvcS21lFEY3nsITuVy
n4P6lMD/WXn938y6rYnnhyCM9CHFlgIxp+9OWSASzpaR+IDt/lukgeQY6es8JoZO
ldzn2aICzwWmLtIB5/LAEWHK4bUoRNhcUAssrYrcNSQGp7ocnhz6lwkuglToSRWa
W/tgHPqsy/Jb01+F0X1nSZLlkVRF1PzeksHFMYgs//Myb7DQ6HtvkGle60fdbrJL
TRwZKrAeLBUPKtIKo/DOMMczG/ExzZLBwBPhl9+Evtk0J7n4n69EVmIPfFPNne6l
ZBAguVP255/zWrog5Az/8IozVnTsloSRtLp+EU9AHiy9cyZ8SQXrSVuDVEDlsJ4K
NVCWhr6Q2K1+zmIF1tEbHmQBincdarid+vjK7/6tpeXu0r7oOTsIwY0lhdYOTnZw
U6EA9WZ3P/kaHCnDYK4D9+V6PiD2tZx+Ym6QHr1l2Ex1/wQ6JaPqCtG40RZpPM9w
q6eNfpNjhFSN2tzVzvtGVgioAmgHb179zHuDe7byaRP+Czgva4YzNgEvHrS89wqB
CyqWXSFj5Q5e/nvbA9cpUdbPgByC/SfFcB9r/BslClpJrgKP7g6649CZmyW2J95v
tQRaZOGwNFO4NJA5/yr5+QjrzzE1MdPvXPUuSL9OJEs/2doNXuJC2pCeaL65rYhm
KOCFxmaIpsniPticu87J6PGwIgd+cmQ8fAnb95EzzOdSvRa19kyXnF3dN9sya98Q
iIMnSQbUaET28qiR09WBohWi3GVCL6C+mrOHqwzsbaGrXUXAX58AyrzFhZmTytOi
xoIwFGFwQEwnTgGKEpPRrW6x2rmkqWFX5Nu+vbYX+I+t17lfQnm+RhRmMTbyOGV/
GqKRRFWwzbTDqHitFfuXuSQ0EZuS5pa3thYjftdQ5X2QEymzpKR4U7lg8u6/bhiT
X4PZyU1tvLKc945cJXGIxOG6g5vkZhBKudyisM4XJ+BDh7voVAraZmGPDnMiUX5J
uItA3LP9iOPiO4NhccH4j7Ge9XU+LYBRY8y3HslZn9DH+iK9+MlVyMgjYz2sCTEZ
mm5qsEUD2idBhb8yQa4IzPFwZzrCLJcm0A0dTOYLcRw1Aq4gTOzxeffh1KxSPI24
SEmt44gpqXEdSk/CBkUvQBqOTd0G0kZb6VCjzcWwDzzZy9fazduqEm5SNillwZq/
8zQeHCj/8NkvIO06w07XTQrn3G6EA2RY16V5Ov5NJh6UvzZun2vL/9fL6I/YsFA9
Pj0HMHYMTvj+g59hvXFJx5lwgCYkjD51Vrg3DUsBuje6L5C4N9qKD9ESJmGFIixG
OHhGUl+2YntevqMzhOotxrhlkv0Yt3AsXiy7mxQgPgAW6diY8KBa2gg5nTNQ4WZW
BZh3p/oFFAOlv9Lk9FBqSSrbhF0bHxDLOiJNuKWxccN/Y+HN5zw99Pc8UOsXa7RQ
YD/ZTwQ9uuaohY2j8tRT3EwxPnpG3UH0DKkMTzY81Ht3/RN29aVvBoyoFi45fevw
/FTGMQpoD6ZXyhSH2V18+d7edXvgNeXHBjuP1r/2wyVEwl+GspCQPhxBeRihUuui
y1ikikgQYcA1WnyVNUHxm6bMspQ1R30PnJBEWFGI3XFUJkydlW/SQTOaL4MS1JQG
UhUFoPFltIHB1JjxoIj2f7FqPQYIgftAGxisSG0G5kuq1N3ebAgE8X8CCu42b0+Z
/pnk4zBXAr03OabA90t6y/jT8C69W+A8Fnp6K/qsz4kKwfMs9hSgv9Qt7S2h8eIt
5xBJ70t2LkkfW+2v2wKGd4EAk297ve1Vnnxo3C6A90Bxqq6AxMhteRYh9JGKQ0KI
i6u7iKK1szb9x5RBTJBS/CsNFm/avKhg7cwAI78Hn/pZQGtfBG+eT1SuTEn/oAyi
Mks3Fm16wRfGBAdqgLumVYdodBO6BjmskR/ErXZs3XWOaaiJgWGiLMbNpOZD02IR
WgGt3APTK31eJVgWYCbsKjaAvV8bsduN2G6UNTqu6LW9BTTsT242grbIHHIv/P9K
4Db3OeXd/Q754g7VjtFFW9pK2SJB6sfELolFNnaCeC7WrrcJcOuCJfl2TLV8pJgc
Kl0nnHIhP+k4KBMNg5FNVUpUB7/qZDL6lrNtG35yzSLDKB+TPcxXGQqSrUK59xhO
w0bqfFIv3N1JacvjfecEWBCTrwaB0SlzY3LtCvq4TK1srCU+zUnjuHNxF2hV2m7N
t55Ekv0TniegVGfxvzzFIddLQNKj6fxE8U+KtCDOGR9jg/Fz5QCpBY/B+MIgkjVu
4N3h1vexrJtf9dfX4kcvvP69ak9wOiDRVZsRnQDcbmWmVRTi2R9WaUWPN2IyBWTt
mswqBVaYmYyglzThWfiHUuS60WI+sD7wQ+DKjMyoLQQkVz0cOoi9EuU4cyCjVOa4
Cdsux3fJMDMny23gKAi1FUM+osxHmU4eSQ9S6B4mCUOFOOXs7N/YQyX8RoSje9Xb
msU8Ao6oZaV74T2oXj0gRoJbQ3/ljXhPfxE0voZPlqKbSwQPEcATEh9v90EXdwtj
NFgxvJyMtB5U25ERBfEIiXA1uuHHvt9y2FoMiJe9dCRpH8fs26/aZ/vETQWv3+IL
5ICtj0LUTpo8R/K8Kqjw/YElI3XWLBa227y+6QkKE9NdiipzqphYfSAWcl3fS48M
9j3oY62GzUFLEoZdnRrc0BD32Q/sqnulQPa/Wd8AVOSsI2gnAqvsO0yIAD1+wXxe
5DSpRErkfyrzHR1JrC15zEQBzx98M27qpkzQ9/jC3114Lfvc8RjQr9In+H0HvLn3
MaJr+7zF1/owy7dRQ/R3lHdeOFFVi6YBKJFFUvOdFgw/YMiPKJUngGeaD7yJSd80
9fQhd26IBhU7U5k/msGVs2BwbHkiHUv548rCWYisITpSEGXP9nYAo1NrnhW4e6jw
xl55kyybwsb+k1k9r7cLpxni0mP9ocLwtlQO+cORbZD8ZadhTPd1yGJx7c431khX
SHrUFfVqZFWi3xAGcdflODa7RcmS7oAu8CB0ovdmWBB5I2fRw1xFPu48rKDpUEtk
uZx1lFYsQd57DyIQGgDPmJn5FmIVeDVOKyXRJy+KTsxX2Mxo+RwUxc8DZACdqrCs
CYAoSrixBSOnL3GMaDeYPb3/WIs/D85LMiFjuh8nJ4WEAGjMHTZrGjTHVKt/fYvH
6up62PQ9K4rxfhZlQjVQ3Y3yVAzTkHL7xfnR/EPgusdtzfRepo3sfYLyItRbd2/P
dvH6UJnmZAJnJcVbR53dRt0fPvikSbk1iUHWf3coRpMB715Sjy/8Dqd14UBj7p4c
XfjPXW0N2hHEXBtOvXT8INAp6+QPe5JpUH/owZt7OzEP82E20V9tdpaGpf8j7pMO
YstVxpaolwoAU9hwXOxr1aNE1ebtzEI5tO5mX9E42exzA1Bf1Z9U8jTlc130LpVy
JbtYJncTH7iLMEWY4UIJIY0ca7ARnmfahiurW4MT+8EnUsAT+odb7hR0PyA2XgiS
4rx1kLNVLWUwS1vElViHQ36i/QSBhDijJeHu49oEwVuCYZi3QrFPI2h756yraOeX
XYo1t512gKTDBve843C0IftLMpr51MH/jlzdsWZUqFLWmIUscLiHqVzDzEbhe1W/
JHP0+f6QTFta2HEI/0OpzJrUZh8y6eudBf3WPTQNIJg3hqLWje56jA1cpBhAd2jb
pivCG1rWkPJyolnbd3Jme0In+ZnJ/2Ytiz6pbXWMabpP6BWaDGGJFAVsjau5cQ1r
MCCtKDWD/w6OIMKYTat/37VlugfWFwyfy4M9c+heVCCJR+VgT9c5dX4LhernYQVP
OZS8sfcXBTlOftnE5TKGHrkrr5SLazQv9ZET8DWz2Jr+zEr13ucdEwNqZptJRoKq
GDopTLoUApdwU9o4oHDriGqBwZEZxZVBhk/nFWNnz2nR3NuQXTznKWrjQVdio+Mb
X5q1M1+MW0mR1fa+iLFUZLRO9A6GVmG4JuOr2YlS/sVDhBF9deyfLlImBpMpcQFw
+VOmCsoRgsHS+QhVLTTHXqwn8fH7b1abibIU4f/asN7DD+PJhMywlBXXlshWmxZZ
W00PlGFPyM4Q6xknxzYvbjvXCtnJ/7R6UR4SLxbqR7V/nr9USHq52glkmj7YPEf8
CLPQ+qQH1vuv5rzHczEpA0Bm7Cc8jRUVKIlA/gYTx3HnQpWdscuH0o0xbXtAZiBW
w7j80PVpCm2vvMOzyCQMO72+fFJ3uMpNUEHBAUCA0xdHm/E5PnwjTp+6THsEPUlP
zrNa4edIaizPPxsXMUC13oXK18YSlb8CqPEc7C3MLKZycfDaLSB1Je8OOIA6D7xZ
Q7Nl0kuEsFQ00KeMwZq1AdWMzkLru8OTVztV1ES0ACJsu8s8DoJL29/5jjpvX2S3
GIEqtm/tMCWoKR8vfvib756WvJHDftsUylpnKVvtx8TiMQs18teWdYQvcpW/ZCuT
6sfV0y1VD/nKPoKASMwvJAbo1TaTIPEnsuWjAV9sxwp4ezmtWo+opJgIVBMJmveu
P4lygTx1jPxXPjD/duREiEghYb30VKW9kgIKdzJFiaJXHbBwOR1AQPPlm/1uzPKU
C1bogJ5QoHtP28UHRhVKmANoEJhx7oETDWaTy1QpwmPd01bszCv/fVUcpDSYbOvw
6X7PAnF8aUnD3hbo4ODIkWHQiOZqSDGmziFM+fiHKI1TGW/DJSnwpK+Mo8eDADO+
34K4JJUCO3SZgmDuhSB3QUJvPUGiEHUdwdvfq1mFKDk/m4KXgLs8QB30O2trLtMj
9eU6u0uIt2EbPrqSE8iRrd6j/Y9rQ+22kPXsswyozB3UsnR2ivmoO/pR+1nXL3SZ
IgTd8uEXlGF6yjnM8jaLXwSSHK/itvfibyEY5w2LUyw/Y9SSvje2gJsZoZL8bhVP
uFF7K688Oxbb+trRTmUCnBE/UCvoahsPkFU+NIEmcS5mqauno2qTyQHwhxW1vDhL
4md2HYxGc+tHzYgJD9Er7tzJ0RBU0TMMxVvXkYLFYni1zeEeOAPJAAE4UQftepk3
LJgHeLNrw6NHGSy/W/srWcYt80kysqQVyjJMD50BBBAzEtAupq2dnq63hZ00zPKY
y3SWhUZyKRgmSfARgHSsbrQ1A7vHjmtc2iqglexqSB678rpYoCSsylyD4uVN30xm
n59HpqaRCnHpUHC6YlAxQujpQ8YQsnkJFHi7AeNy6eBWdu50p+X/hLU/HKXzNvxh
4OMf4teSKranjHYQs4UCyDgp/MAdt/ygfSA7lzo5CYwSku2hxiv8hSq8n6/HiplQ
3+wkTLV+D9P8radYUi8TTwvDtNnsXCpATRNqwceg3jqbMtriDsyan/AbDID/gcF+
H8Y3gZ08lfOeHIXhzKg3UysSHBtjRPGXJfAjxjuW+e/RfCAo7yYPj5vH0kNT2xBJ
k/lIGLeMT2KTBikHN8K2bB6dke6aHn94+9GSQNhVUrEgFr031XCPiPVi6WDTAN4c
EOROig8RLt76KMg5ndfmAS+zL2lxWtSotdLw4IzQSObBqvg2+efkc/8arBG5I6DY
7Imt9h25z2dwZLi8s/2XEDSEOiF24gbSdc9apQPUVd7UrLkNQEXbTZLg/Cls+0XM
yotsKIxrZZL6e3mzkb6qopE0gg/GJaiQFyejIHKt19A7pXTNoR2oMGR4l8Eoeji1
CdpNTBmFlmDq8uV7l8/aSNSqcCZVpJV0UwAabxNewrsjGuXDGQ7iNTwdr56j8FdB
AsAmIUwOz/pQCWo1wAnWSKVI2nm7xUvHstc0jbt4gsXaIdlKYLzJo71T7PgukRKf
38QfIJ+HYbozEYZ0AQjVKFXfdza85KgFnFiF+9PzqLDdeTODfAp6Fr4f8LHnmzAU
D2xLSlUKkl+lSSP3eFA0vhW6mhXiKqepYiDwlwlQhN/0RjSgxpYefUDF6crfL/G6
jqTu+N1USuhpbAmJv4PcZ7xfRzxb9Ga4wbwcPLT/plNt0kppN0wydQAnjuCq/g1x
RG60x68mixcD/mpMuYgH5OY8562jw/oiVn3BbmPGPljYolP/o3C0hHH8gK8VlP1s
WcdQhe9MpogOAnTSkK+tvNENLltNJeQ65vWFPvlas6uCpOa7c3bDGbYXdK8JqWSh
9+c+LfD8g/8Gc2JYgLcmvqB17R2b9Ktbk3qvVUhTbtIig2FW2+3BflghhV9zy9EI
zeI78/IxKd/XvtcPDPr5nLOkmALbF7h9qjpqIHAr7dLAsOCMf3/LU46U/BE0fra9
biFI7YIdRLADBaEGGpRkZkAJ4P40JrpJaQo1ozINmIfcDdDf248woDfz3UveIopE
bhZ16yr2NtxcHxTSjVVsvAJft4Ewtd29pf1cxLZhBQ1dB2YwfL7sQQHrow8lXk4r
KKVQYwBxb5Q6h2ktSg/X9W+11/iDWnxZziehysvufSvgqJGTWbeEzv0yAxF9euJn
zUWULBkH9zoCnHC5GSLj1F9pavXEpxg5NyM1reI2IoX3AQ5vyJVqMPy9ddZv3pFy
WKONVQkW0zMsegDjtKcEXt3ZWJfJiNcO9lBC62qYz9I624XCyg/oxsRiiKmpfJLQ
AG44/Ujgx+NK3dy7uj7Rp4viQJCXtgBm3LK1YHfaoAHXD2y9Lrdwk2UVfY8Gwe+7
MN7L9fzyffqWzTKeDxgmsf2eZwkaZuIWESGcX5Shf9WZ0o9vsz2KolDOxMXwtJWl
mFAg8SbjmluEjeJ+LvtOtjpuRsvi2WPtWU9CpCAZI41ySXQi7R5E2rfYyIpXs/Ud
cno4vagb58jBsnQwK6xE3EQP0BqkWOanvW7yNLdWi2cyd1SATsjfwSzMSUxpRgV5
P0nmVzGsimui9TcH3yOuWA1pWLuv8Gt6OeL3PGGtlPPszVwThqZh4t9Buhn1WSRQ
UhWGVGEjvU1l73o6vfC+B6QyVe59r7dotWT4EwLycgz30C8vUukNlGJRWPRXLLuD
esuC0ul2pOnoUst4f8GMaDH/gIoKNv+0us0tL/StGD64IR+oBlodFf2hghO2tdoL
Vzzdf4T6qvso2BYwbaGmzv6fshtx9gLm/yyVPNwTUS/k2gEVMJZZlI/LGvrO15yq
0L3ro82YfEj+/iOcJzrXuEfrYmbPvdOMSuuKMWEiFCBaTCAbOG+D4JL9X1or9q7g
WiIeAPzNtpTc2l8gnXBz5vtUmNsbR/GQePEFR6VzQmBVeWMs59cHH0NannDEWF4I
j5yWJWy2HPdkLNrBOemo9Kq8ReJJE/jPLIz30NqNpLG1fez789F6Tz8zKMg9qS5t
Ud6UuEXpyEblnvJAGBJGIhZyUuFQ4s4zPlPG1o5M/0H1rs+wLM625TEFSynrBA3R
9DhU9Po+KECImpKSc4Ra8esMG31zw7E+iuWo1nIEkhyR4i3Jvz+6BpT9XJVCjTgi
hhv6dLiUmadKqc1Q/b5FjFVq56omlhK910aMwWg/Y6hsGMqFovcnFkr5LgJLWjFa
CPUlFw/kJX2LddGsEn8sfJdpi4drxk1szt1KecWoW1ppWdpyIatx0bQVVqikDaGk
sFuYP/sMIABmdX91HBiypyFMZuRIg8+GhwZyjt9H35My6M+laBn5mEkG+DXHYA5s
1KVPA5E8CZSELgnjM7boLfdGWzo8+Fq+LD+5CjFC1Qggr5+HFa6qhLSRnUeFG7ca
+zUKo15LTBvDMUKtqFTZQXuAFB+K3FOsQTLl2+vnY9jjpyqfgj4H6uc9sdqrC8Bp
uGBZff1njkd1Z2WU8GlPV5AfIWDe0D3w270MI1ua0o46BhLPZYeg6RimszdH8Muf
H5qBkTJVFLwF3hwp6QsfNtksFzrRD4IaWDq5CjDcOfrSSTa1yprWIWw+ldyBaWTW
b1u+PZTUIX03wO5B5Gbs2ixuasUSTpjklhlsojWyMyWFR1RA5Y6DJHmNalFkSiiQ
w9ZlqWVfkJBvjm3YaUJuFLN4vLHzAgy5XL2hQy87S4pyP3pXFMbnRArNujPkfLas
5bV7MroI7/VYwOObjSjXigqilsBV2WE0DZCG1rRqXz0MNMX2csGKPkfT1Wfg/rO8
AQOo/p9APYQSZjU03uSY/IyNoYbZ8zu0wd8YU+yh9BgALQfB7TjriruYeVc8d9+T
QePJ5pO67pPphvpfIWoKWT4zrZK8hfxa07ir6g2NXHzOBZwsZaXgsymr2qH30XWR
rDQ+8GmZDnb4/YtHIH8FOsAePhKdV6fjUUjinwSxM/49tdEi8M739ndGnV4RvJGA
SqOMAY3iCSWnzSVO7ytlSPdv8WLe1tw8qvkMUiRlkxz5/CaC8/nS3baBFGmzpH8O
ELp+sgE0XDfyhpYr9eW3kGMwre31x53E9V0TvsbCmMrAVQuoXSkW2/fV26RLLQ0k
1J9tj0KdZlVlYo55vtg6UowvC/PjHb9eAt3mGbNdJZLGJ/Ee5SaMJ3xVe9/ofb6h
4su6BFtxIxruxurv7RmsQEMp0MpDkhz5JYsGEAncqTzKtwG5ADmBDSU1BHvmYR5U
eG2HpW5pW1HR76uSYJnJQhxnGe5u7QhTs0SiSyJlqlzPrzig3Pu/dRukgOD2xjQ1
cdzLo9urlt2SyJs2ksxGTPW+Yak9BSvAGt4bE0aUkyu17yMCRO4FycNiN9fKp4U0
jBC6/wEJF6mVsLcfzKS5eS0Qh2jM2Iz2Ad2PMDuGykSuobrYOaMpKXVowRZw+Ai1
2/iIQ2DVTylsOjxsa3Sh7oy511ncRvmPcElNIdYgkwG9NmksBZy2rZqpkTMbqOgk
9K+V+SkWV6SwIJgDnijHepbuXCWF0VFzafoVDZoTGEjIBLdFwseLN4g56mGs43lt
7IGjSQE9E35+C57jYI+USH4Kycsln+54ut+LdqqyzZSCBHGmchUdgECbP1v13ChM
8rG1QrM79yxJSASJAZfEJcxF8n1bNOeQMnrXbx5fMrJwKq78mGB/xqi7t+kTloqL
gclP8g7vCunujCZ5njiyDOSksSQYgwOs21I/mxX5+b/3qICYDIoV/unm4wONKkU1
rCZieq07WrqRDzrTazYFIVE6I8A0tmnenr62jQM2Yrzv+917PC5wApVdpSrgdIed
mGBOkaU6AldmuHSJbTZ7qsR8hkwiU0M1YT44XCbnEFhZ3D0bGDVwnUKWoGQl22ze
xXju1VzdLRkqbNyNRSO+bGg5+dT1mitOL2wcVH5jRZ88jyea0p5NNQAorM1dWEAD
tKwiwY4azD5Vg3Mu8Y1rGwUR8Gfq7qMEQ880RiWdJfRWMmgxT6hjW61jIOpKbCyq
+MQwOaMKn0sHsYY7nc8lfrfN5A595hRTsxdanwB5eUn6QvsmBHc60zNh0K7/8tbE
F4CnJbriHMCaRU9A/inZjv+NQFz0oBcwYCiKqIyTqakp4zs1v6PIsXZMBW5dQTXC
Q+1JfMNunibzc9qeWl/cikRXFIOSB4j/3sNHpZAic7TF5/zacAnBPV8g/lKXb4O2
M7/2QGSAK7ruqCJEHDJFVmczk/rHj11zdFfB6gyS6qUDDirT261WX5irG1skRfGg
n8jdR0FWdDHPArrJlEiaJL5zOiTCUPh5vhSPsMO9RmeUdJnf/I/bE1Xfpj4J5a0n
nCs95tPZ0ceFY08O9ZAvA+8VEYsYbU3gQzb+FYjQgujE/2NaMaUOBT1o/y1qMA/I
Ph3ec6N1ln2UGlbzNYwWIRPXIzhS44j+Og4KVOFfYmnugJkRVyW2nLA21CmdAjhB
8ZIqHW+VKLUEob1226zXVf1xnRkIESFOerpIYofGobPL6R+8RijCRXJJtcmybf2N
q/VVaS/ydp92izHXag/RqyRIJ6SobJIUg4wcp4ankWlw6wY4NXOaBohRQWuIUkTf
W0ToIwmfYHnph8PPZEfO6nIo/g41MYcgdKnjJsH7ISt65AHM7bbdDv3O3LzjoNNC
iiEwJgvarTwW2pzqJMX7aO7G0bo8jPN5DQiVLd8/XMiyoVwT+ZdqO1UFCvsxLXfQ
Vfvn+shEQTFhaZuxCd0p6RIaVfNLbkX7DJL/sKhkGxfBklFMEse3uCrNBypIXCK4
9W7n+V0STeTV0HN8n86Zvshg7a1yredku7FeUIXYD0Frse0BNnkLVhalRGg8BxUz
IG2Qc0jhLCLzF7TFGVZSqHf5ClGSZcFK/Mb53qVicu2vl7MvZj9GTZR9K8PzLEsi
LNpFA3In+HEhSiM2vYLxftdwDLtZWG5vKTz0HzViou/WB6aZIl0w5M254mQmzU/F
L+yb2BwLC9u5HKWp674rs7Gt/13ynUa4K1MLpdT0yZNKqAvHFgxytg7Ix6PhFG89
tVsepUX81TfShKLxaDoM1rIYS6qhv1lbIxy4hCG6H1xFJd4wMC1oEV7rbfqQ0cvM
EMEBux0x/NHoTBvWQU4+CfDPPNe4NttF30PsEnYlqYn8T6P6FRLrMziPRnGBIkEP
58LaiUQxVhWmBnCPo1L3wyczmF7uzTty/bpgoet6Ya2ui7/2pu4C0tVEW/TOtSCG
UHdKC+jqvnweSZ8X4sJb2prvCq/4tHfXzZ0GxNwPfLaUfaOlsgAz4U2ujrhGiT2v
B6tt/aNdD3/8hAxxwtWxeWqf20cF+XgqSxw8w66NRiVQTBa2FCd4kTZSu3bqTOmN
bsZdo2VmNBUusmmS3ER3LEAqWtiInu8bX0bMxngHSiP+KrFw9P2SSiUBE9wnDQY3
uWvsUzNEmoTrDSZTOZ78Mbg7KrPsZ4Yu/n8XOUpqnnA7fQRHD50wloe/nIv/6TY2
2Gtvq17dj+DST3zDH7+2wha0B/r8jQFPd3DzLp1k5DKreFDxMQym4CkYgb1KDpM8
ia7ENP015ZPwJOBjtcLusjpaOzr4D1KE8yDgr8uyN+PzK2gMSonZLpe4cuEAe01O
yiJ+CoR5R/nTv7fx3VZoOyWTP+9qZPHG231ZPtq0QkLNOEWpoX20ujG19dj9pcOB
Z+c5hGpDTVz7dPYAX5c4az6JqzhTlOFA7TPQ9f/iJMz5d5JeZCzoCJ0MT7YGqjBk
ULr5mSIfJ7zY/wTYVAPyMtBx1+JpHisp59sPYOShxdtwljwRM6XCplMkmZNNi1GQ
Hqhr7d2ztH9u7fzSqUeVdyekxoit754++GEymQGCP88W4btWKWX1DSwYmUhGm6J0
9kuK5Bc0ibwgnJFxRuGolmw/zkwDQrAeYguJLXTLFxCNxDt5tRQq4bn5W+b133AJ
5K7GGa6op6wMMlpBxYLpr6mYNOUSOci54YmQCVJRWN9xR8+pmziKPe9YEqtFAlcq
FNjwcK1SGukZ70wRIpb3D9X/a8RNYHXu8MIftMG8dFZBrWNO2lDUn5aYkCV1YYcM
DyA2xQ4jUaUoYEHLJGFP/CdV6h5XwOsL7M+zWgOfwpM6yXl4O2qTXydaJCVLJamW
T1dfL7ulcMQC12UqpJMLuRZG6GO4192sFoljtHJDJ6S/lCd9QeZuIfKEzMcCYNfk
mb3Z/Vex/iRBn5A9C+ggHlElY7BORC6/26B7yYsELNKQO5GbiSYOLVC4DOekj+cP
4WQA1nSxcHSpnffoIkNi7tOJyAtG/IknsOopqm5RRVUgOEMSBmspT28vE7QalGS4
vhc7s+V6nHLCiPa8w0PofXIdQFe7klcD6d/5AhtzCIDwJiPVyg+XXKGjJXuJB4/Q
hzoITaj3ypajZpDIEK3dEaw7/B3Bd6z3wtjFt8+qxWgG19eLZgfpcHQcUqUjQ9+o
RMvDDBFIn0/Izv21mFeo+wRBsKdRk2ZY7UKoEvOoydYD/FOHn9a1qW+aQCkYrpPt
GloOxHkCLkiqHubHcXoCgNx2Qfnqy8ogtgSoLfjajtiXrTEacSjnsmvAoCR0qYLD
pgt3ZbKj9U63X/9CH+SmjPuu+6KiKiDk8/IXwjbucd/acyYe4VbV7EhaoHhlvfAV
pGiQBG/LZr86i+MpnsSXHvON86TjIIKB9A1InE+MLpaI/8j+7GVPbNx/2JIt/d1i
sZWF5IsZKKhhX3mqSTqeFZuqq6e9OPkKcOVjrU9Q8IISwt3NUbP57ZZVZiobCdhj
AYa1xMjGuMvZS0ywAhDgBYAHXAttzTN8YRonNfQDSRrz14gNy8CKzQjsut4xQyBG
n5inArCnq6d8EUKzH2/xvWrKs6qky0nvUzO0MPk+/f7qGrofzPiaqvKrhcH34fwB
gn9HS6QKJbT+RcNQ1d9TH0F0Ro0PhLQtkcCDIxdiY+FAH4WUIPb/SgX/4lI2gOEU
Gia3uoEqr9TbLonCxzyEulND6jJNnyXh5IqDK7HbEdEkWIep8r6vmOLpRYW8fSHv
emgFH7k9EOKIIhy2XBCFsUyVVT0B6AU+S0/bT+pW7GJ5SxVVpbJRRO+vDNZEOblM
3XrE34ycmVlY1woNR0GZih88M0+LG8FBD8GJMF2IVnsnnlteR3WNouEI8mgUgCJL
49Lzw2FEjPj+ZEmVKkmjEnq8l1cQOhvHpfhqgpt4EMjCF5pOX0VUkjCE9jMjLPdA
W8mg3YeQpnud/ZJE3w2oc/OIqW8NPl7CVEWnt83nhOXqQeKq33PdmcYHKHPGN/WR
IIqziQwiSbdAAIVHg7WgTnFrHjvPhFXhcomNGN31+5yDorfsvOW7upvSrVVt3vY0
Yqgt+GTpH8qPwdoZH3KSx8nhGLhyZw33ZAoI8P6BF07v1YF19jf3Oa7zQr/SWoRk
nZUaezaDSV7HarJJ2kO2i69pzir+7P2PfciwwOMi/Xc5IZnxtXR6FxhFdmJSqrOb
bEodLkY7OsUms0gypaImWdJRyhz2qcNVtKR3zA/wrXgYoDRs1qaej7Q++UD5n9lR
3w/xQK99fwpqy8tzDXxhGm+ciIO2yN5k8e5g1xaVptD9ex6YSnLc9S1hqq61in8e
P4nbfkTfAYqXlbGXhD/DyjRoBs+EHgHLsnoaZJpU1ruXtDJEuP+zcOb2wo5lOpxJ
5EK4G47tmjOYgCo/xBDcUyCS4UkXh/z741go3sLaJHT5q4nECMOWNs2leEt+VGhH
NbgT6G/De+iT+Le8gRp91REBb9oLd9dyiq5YBsmdM0Gp4DP0uBddIJJexPy29pMz
7APBWTitnCCGd6CrOdl002+4/mlOPltT6tZz4cV8NSrl+maaBXtC1rukebaPCttc
lZFBdT3uBQHUk/zH395D34j5pJqH8CbXwHoFFMcyoxXXyDHUqQ7uWXMovJjjHtUa
p+rYPBoeBcdW129KpUUuT0zncq6knxnAW8NeyVGTg5RL/KXIm1w8NlGQLfuuYFRk
VMnXSG8a2YkBeFB2IuLp/j5IH42qOrCQnPWPlLVd+Lgh8Je3JPJgw/gFu6Rm60qr
+KgZ/dVpwEAYpVXugJw61uv465XtEMU6PdPAONiVjQTH/s2QOa7hj2wTGrcH+GfL
DFKmg5B2YWoU/CXDcLsGj3JsA5pRg5SeqKb3ZHthaXVft65T9+gK++5dIVj9l9cN
t8CIRHzEspJf380pox3UTzcTVmKvXBEAD/xWg8WbaqYGyyJkafwtaTnMzBWZNhov
FBmXjwPiGh3w40xkS2uy69C0OFRsVj93bJNJjB9tG+XMsfew/fIdSRrmUAWwoqJi
TsUjyyA4IyDaFVF7bdIrzO5LSLHl6lhJiLBh6CmlSTCvu1YtF8swhhmPCAnxK4sM
cEb8vgUCupgLO4NFYJ2HYCv36Yxzgmj8PtJn2zafwzesksyoUzF4LDOVv7zQFpOx
PwbHCWnYU46phDarw61VO8apTRegQZXrGZ5Is9CnQ12SSGk9EE/8FEP7y650pANc
B2n2pXAtldU+vqAEgeIYCASCOJlVkTlCXgUqGkBV2ck36tspXKa6aqBLupOw419s
Duxf00MNJ3/UPtJgiWbPQl02M6m3oUWVaL1+Ujz8chqg7BFiceDmyimtl2kNQRMr
bmBNilZ2zO0ZeYRVZrSI/wuBKjhBADflJw5pAoXRwVI+0tpixfhVWL7i1lbjLTwQ
Rqx0sWtrIGWSzhg+02Uf7M3kubCHmlxb/QVzvCizhTpjOpOeLzKqG5Z4YRgQ++CN
0aqj140vaxmBKX3uS2t1nBHfY6yez23qx6jm+qLiGlcRyDkwTt4GV72wWLVAphp0
lPUsbCkmkH6y4Mpt3Cyrmrfihbi3dTjDMYTFcCyOjHhk/D1adx7IxbfLxuRfpcNF
HkKq4MlBr2W+SStxszUeH2NLCfZsyqzvljBCLIljCOcfWaKw8wOydPdI9JtHrNBE
eiJNn461FZ/zhYy8M6e9L/mz8mkcrQyfLvh0Wc1MX1JD2UJXFpMSor6G7u18YY97
C6ZLGjSMnuHSNGNh80X58vLfHx2VV8f09e8FvFD2XRu5npI3Eb4lo/9XkdzVioyA
yYDk01w4as5soyRyQYBooNO/zC+6HbR1oEbbF2faZH8pvZlypn/9Vaidu+RIZy1r
cgeZoVll+S1/kiWfemD/1bu7OcWPqt1qUav/3tVaTQRFLz4N/PX7MVJfKEQDo1O6
ACD5CN/eRsFy0iqzqud9G7c7Yh+qCar4XU5ypTCM+Zsol0ApCSYSRs93OIV6Xyys
mrt7opNnCx4OWbpNgCXhxpzlq4NK7EHHDEJnSNZhKkp/4v8DTUsvNYhgmKLOOjyA
HghyUgqvwjADQLZYxrYxINV9cja7cT2Dcc/6gjl9iJixtp2rG2JkRVqA3UC4YTpS
ux3GmpqYuovnK9qP93Bo2dX9P38fkc35AFqFsZsgSfbfz0YmwQ6Pf2aJ74FO96fm
EzSozmIk9j/RJ/DjBAKhYJPPAW9oHxo5XprMw4R0cOpDzAeYg1VvWsv6GtRUY9/+
qjUa0X8rmryicqf6p3H4r2Kcz2IOPLH9XbT/FmWmaZZ7EMbEKWACceiotxD8oxe6
u9HJAra7R9jCyU6mBsC3q2WwcAf9MKi+J5GP9FRMZP3+/u4iIIYMNiNzsw3A1TO3
ceYKNgu+UEBa8jXMb0Pc7oabsscqGr2JkKakzsLeNybj54tLP3ut05Sd5TcRIe9A
y6/JC9fGPY03fWJXEt87TYgwITamXiW9Mxa8W7GWhlR44k1yJXETeO1h/OxJYfPP
szHfjS0dcomj7Kid/Uus4HYn/OFKTDjprmWBrhkSrN0I+Gq+hdFzOnZ5IX2824NH
4J7LfaKfnW5Ygu2M5UHNVClBoYVxFiRrVDvxUMM8WhvoQWcuBI+cP398KbJEO2rM
PxWNDIOU64pWy75rRhHDmZRnoC8oxjFXLkkjF3f6sbysjCIju+QxDu4iltTenB4j
4qOu6SZUGuSVZncztzwSb7FZ02LUNNpubo+VJujz83ckMgVL/4KfG22x+cDj3qZA
ZJi08LpYdPOKsy3jkvloANEZwgpT8pr7X9DfGzfOpvvtVzFuKpS+avMzMpe7E9Ec
WXDZzf7N1ZbDMJ+AVndY2hhbR9KopdNJhA9XTf3q0vPmIiBEor/+z+yszxn5aVkD
7z35UlRqIR9cBqjR1XhyzjBVxXc0w2nh4NzdjiNAe6tKWpuWh7FePk5xMb21f57+
Ww9VWu7VGEKQCFQor7vgWY6sJqJ5djMD/TUA+meuWVBIy70sKBcndaOQ/ia318rA
vH9kOa1PR7MM4RHAcjceoL0qOR0WqtiScZR3p5spHyYOQIWWDVovcK8mj30YIwCf
9gAWpoAWVo3GshP4b2OiJGvQnSrzdTs8PRtkUlx5cWnJ15iepBWhJv0sExSASEqs
FSq6Cp9Vikt/29UbzpDg4t/jJk+4vgsstgHLw/YpgiyrQ34BIs5+wxIuXRaiHMcQ
rm9TqOf2kJW7rmLMiCo3uaitFZh7niYm4EJNEkj9UDl4WkL1LuDwmX6x1PCf6sNZ
tgWo9cZ4fWB/x6YwLTECdTWqKNES/12vCKVM0UrUZ25s8oipNjyBT4gNEutigFXk
Ox1KWelf9vHawnNLK+f5LIjGwP8qb0Z3kzlKFoe5cWIv/7DXsCSRq8rlm5Yu4V5U
5r85rXkuFSAstAl5h/vtnDahhFa6pjqrpV6vNyM1w5SxbvON+I3fqLNsygo2wEeP
M+pKA7fqQYGcHNYfzNKyWr2K/WY+tRjSVNY6WUq/GzQwt+Wed0UTz4Ezkluhub1S
DDg2hm0NsI+PMq8RARugE5KmS32lzvFfAp1eifZOKX8mkZpAaxSrZz6uQWPU8DO3
g/W1h/hn/SGvGEVQ8d2tTHVVHif5Q8Q2/5fontvdewKCeoOCiEc5YKH1yFFQZERS
moV4OP9RP0nZzjXj/obHCA5Kw8KkLq0PitNc4QVIQV5xBvtiIAMYyn5ZftFa2Sm8
9XnDjUz2HgTqBTdIIcg9j409kDoCmV1KYzvyYnBSpNPlwzA2x+VBkwGkOaLe57Ov
+oeG66i6gBO4rKWGUOZx4uoGXZO30prBCJGJ5OnXnXCx7JIGfO7sAlQfmVU9Z5B5
6ZlDbMaSwRNlULVmPmL5k9kyjEP/31Ez5oIsy+HHyGjo0vcNZEZ/P7gv8t+VEBus
SctKUpZzB3K+ZocmanLk1I06nxNouk6kA5AucLB+NeFzV5KiBeXDbgYjfOsaqhG+
SMfDPN23CZv6B6Sw7+dVrxza7I2eIfyBh2CqT4wYBeFy8tSnVLMbB9UaQmJQ5x1Z
ElVthTt9DNOW+FyLv0e1BBfSxdMdWrnymb4z/jM31C+i4ecrUmCHB/P2+FAUH6CI
GtICjCu7veBz2RUgRokGI9Ug+0Pf157Lv6E91F030eLWYvVrF4b6I51l/YOw+/af
30Du/couFe4/dT5QomRdRJCnktrfnlzyQpDb1yRo6csAT5hW2ee6W+OGT38sm19b
brsVLvcJszaj+Af69l3CaFURsxzSh/mUSfecgJ4lQNJIxbUB5qz7tKgl4niLWHHP
NbFaeLOVbeJVm0QbK4x7+NDzgUL6TbndIRwdEvQOlid+qzVfwRAfpwsHm33U/Z1a
o49yU2qLMd5ia9NVfV2sN07hfqycBRcfJDvQE51C5Sj6c1NnsDftFg28lb68esf9
TZjxX928vjJInjlnH7AJkJXJHihmZbX1/+bx6mGVt6GqDgZ5hbM09TLlV1ST5ZZa
QAdZuWQ0x6k8Pm8X8XWDQlGye+6ljhxDZS5sUip3kG1juoBoeZDJvj4CVsZaSBRK
wA718gpnOT6X2fM7MIVQ0Ol/nsQ8kimVBEvGzLDW7Vk+NT3NoCTNwWB4sgD8bCvJ
CmlQ9NwNNaHnmiBpvVkS2FIkH9VByS341IuZ0uwc9UFsPd/ae+Q95m0gKXwa5+kf
Wd5HCgwDu/SQ5IknXMJnv65cto4BDle6keTsA1hCiw6msklFY6c2HVTYrcZ19sqN
hW9q6mggDWJNshyTZ1M6wk0M50NInyxV4sVZND8H9Hn3uiyaOdq8++n0KxLYLKl5
mM0HNJ5kyffFw6n47fMciJ9pbzu0m1AAP3jvNnaY3Z4LunKnSALE7aIsHtA3P17f
1+n4Il4JwaajaYcO7U8kd6gvQW5RzRMSWWyTCizQ7pTLx3OOqyR9H4a2mzOeg0uA
LvA45r/udsfG22KO4M64h/sJqpg3s6NU/7NgrEuOuVgvPZ/Kh174F0XgWPaWyxoX
FFLGy871JBKb6Blr8Ws8NFo3J8ojN9nob5FA47EBQKkvqwx6CfNRCmXm9eqKwlWG
LI+yyp0bGxzHdyeTUDUttuvnGwzJSPcACrgH4T+9hZfhX6ORrttNULoKJ3E9coAC
P55bGtDi1/UDicjQmTKSbP5m6JciWcvYVeeAm4CV6bzM+rcMjrSn8lXLkrhi/D0B
Atm81zVRAQtnIfnDYJQWqdATzIZ84P32RliCtcUJv6ofWFZZVzGPDTg9ceCx0vUK
wVpG/JIy1yOGLrYIcfsPBtVILnjV+T3M/Q3k8hqvXPXM601sWKZe2ZzSx4AxPGMi
5jwBG14Ga8gK/7wYF88daXHDnFJsIIctQ5MKTReDJuz2/RpvOinkjjLpxq6+nyto
JRGu35x2rA+UPPxfvKATg5BlKdjSf9/slgd/r/zd3NWBXty5CT2OvBqcFy5aaGOm
BbXUH3CFaJqAvm8t+h/7z0u0bAYTUkKGKlZ7aaA5n+rbcvsm9YVK0OpXFu1Sy9gL
fjkvkYsZYEUxZw9/ah1n48YfghP/gfFObsicCVaz24/k/v40h9c5MLse1K+OO/9z
2rih3T8k7c9QAGAz7eQsd2Ryu4EiVbi47BKpIEovCaKrmqoHVnXzFYQxlCiUFnta
i478Gx2DBs4o7DiNJBbD6u25QDDEZJaNvN0+8k/e8qG5C4Shhy2tg27I2Alws3TQ
sIhQjhghRdS3UC8E4NOvDOWOMT4KGdbMlU7d2oldhYa1IyVWvTEmOVsuh2U7rFCw
Mz74PJE69uBNRRtYvfzUrQAOZL1g0uWVGRzUyqSszkNcGx+CLKs1vFxVdMKPdRtW
QYydjyT2SiEzV6pVsMDLciZzNrBalbJHonkHOlMLqN3KV0kEEtkN4yMYk8jIR70B
GoQQkriL0/XAg5DTLJK0sNmGZC0hUgnlQmiX+GrLrahEBmt4ulko2m7p0favVFQp
+YoAkm6prIrTaluPDmo5xkUFUIkL4ERPO7sf4jXkg3QajUuJ8Sdva7walpt+r7WY
cbXxpj1dJu30W75BxWhAf4D/EtL+CC0oqn+8d2bU7vJXEnGEdYFMc3eXRDIT2V0N
MTQn9No6BpRVOzScER3Y3JTJCIpfUKwiYDR0CWvavMo0jUkZuZ+YEKhyoxFUxa5i
OggPR1NiiyGrVJcpEUNePeO22AKududpy8FP8Vm9rgoSiWEojEAnWDgrwvUSTW4c
QfczzLVr+CHgoIAVOFAX/ogrAIDQBek1Ad5z6KQQw1t+V/w39jBG7rJTGnQiITbj
zQZBQygOCdmFEWtM9CPo0QWOB3J+RAVD/y5exq1ihFDv9JV5WpUUsLhZ0L580pLf
WQbvmqWAzEzALoj8uCF7ZipA7KxH6Xo3FdBAspp/a2Z7yOs0hHXY5UIeCQJ3QdzN
9CIhDItrraPSxQsV73xhEjOjdC6igU6IzoxuMmfZrvIqn19MH9tSVoBPQK+D5dWt
j+QaAu8u8U7FK2GdtqpauQVMxmFyuNRQb18niXGht60mTub3Iiilf4P4d+WXHQke
ng9RaDOaKqivOh1fDGVN57tGBRAJduBBk3i5sbPBqWl2o+kIGOo/7rHwULRAeN56
/gxXK+lZQZTEo2zrRnSIhKOe4Hvpvmj7ZmR4HM5GVApkma/CXPt+HWWRyp0HVWrr
8+fVMkr7NBHpaHpfRlGwMDRoS87MCsrtAMdauxxrRkGHtyyhb5fXiW+vjMLPt8l2
3whKZtKkvifhssm2wMcxqbrASwuQlZRv0qzuTU5cuceEVT0xACYloYZXFE/JZ4m4
aXCkkVU/Y6X8mMyANjW78awAXbIv4xbEie/9rkWJmHmnpyVjwi39I1hST/nTc8rz
/kQFUiJ8dmT8pSY+Y+GFz4ZukLZ0qIfZyExjrePHAYCBCpP+iCdd41N1sWCRzcH2
MXLGDc77lCuBrT8X+NTheHJCNLrPgn/cuve8bXE1oWSBhEgj1DvQKGciZ4j8Swso
O0gVUfXIaLXHkaJ4p6/G0ccROKsfgxsWwNQBKMp6vIh16Gn40rL9MnMKfg0l6SjD
TJZw8AsWTiEb0ChdrjZ+7vkJejt7AN6x0ipqkRjPhvQ3TxVPyqngr9RMiECS0U8S
7Zetjt5wizGsLkOLEyu6IaxtXT2I+w3Wy3kG7o5O4jJngn39Id6Vfis3uGyG4zih
S4OPo6fvRt69S36P24MWMqlYn9EJSItYDsjdLI1fIIWtlu+Oqbb+kWx4LBZajXjk
qBsqS2ROFnqTQccrUGJ7vVAPzefFwMyXF2BYBuvbh35ZqEyD00NL8TyJxod9aW+1
5zJ77hMHaxXrEPouNF1avbfJJea3si/vJIlHwLgyUJv7is6V8kBsDokoZXCvLRxH
aipvJE6iMRwWTUuSPt24PVDJ++8fUsB7/46yT/l2/a0AUJabOnpy4QBzOdfRYJRw
fYpMWetSuzluu9YEG4IEolg/sRHzTwvK1/NY+FovKEE14ECqO52lKjEvtGdmJyAR
b/LySCmXTYlDq/jkKEM3eo2lL/eX1q4X0k6wqglt9c4jvhg00G8AlcHzt+seYNNI
qDzgSRNe4ydc9GgCV2S1LL8/H7C4kn4NZlPIl5QnSPp78tM/+OFrQb4wFiRSN6UF
lcg0Afr9rViFLiJQLutrQjdAT5lEnB4hfNFF8CqpVvd4MnuOIMWrU3+XOy6ntthq
ZRxVh1hWpJzHls/NV6sgO9EpX4B3Zvis/0+NlbCF890xDdBX/x+y7Md059vPcZTP
JeUakhVEyamPFxj2pnOhJQ/jCY4n5PPkC3zm9Y8urmYlBhAVPT+fFzyvUv9YVBdL
je6/WqAlJpRH4AtvK9Cn7EfQ7IarN0w9Qill0sFAATS2fkZ1aYa0umxPp1zJTp9u
mNvks5PAZzwF+oW5b9y+JPVdlLTEGe8NI5TQxc6IKHJ4IAI+y/W6blYSxFmrajUP
euBpmDNJ65K9xhJ/3zha21s4tLiZVGnGc7DmNlBjO80o0vmCQyCZxIlivzELeE+z
4qnJ/kY+PMUwudnYd32/0zQ+Va5IFH2jv0VQNg0YLRtafnborjhySiqqki0MBjhz
OQdqjaw3hF4JCvmV52AJp1pXiQhsYq3OEOFJb2aQNK3YwrgckqKhna3J1Bk2/WNe
WVO3GJx49gZVtoinRbmAsfQBnV0qW4PXiYZlIsqrPgH0lrz2ha370BaS0kgaZ96q
AS2qOtEwVSpOqwlNDSyptcUsN1XNC76RLCSNzroFJRrqo/hAMPFt41cddhHzbe9U
2qnc43c6BcXnZHqTR6gQ3vY+7FxWl44Qozg7tulKjO7Lj0QUwvG3kXHSBUCgCqnA
MuN+wUfUI7g7SgbBViDwJp+a7OHr7Ma/+zWaKEN2dfKIepUKu8pE8rdX2R+4e+Hy
tUBX+1IwHKCHHk9htdisIPiefSX7FcZk6B3r4ATdf4qSe/DpbHkM2WJpPUzIuxxx
d8SaUFZjaIgXZ7Fwgme2BjFzKt8KdIUs52Hyfa0yEk2bgb7bgR3RdEvBJVLC2mxP
JchKsN1X0PJx/LOKi3JUv0htUI5/QazW3mtNHILTt5DPdt45ufLjroH9yYcMSx0t
dk1SlSDL9uIIZFYSjVxico4kGiAa88FOSIOLCA4ygTPTGsRUeQSfXBvH79T3eOgA
GKFM3ucP7FAXiG7XB6x7BmADStRsQwNyjP4JKM66sO7NUMoGSw63qORNQJ58orKm
0JY1gOgxSm+Yexb0uAr9opQ0Au6D6pilB9P8PZ4b9ZBeMSJTbMmsNb73QChZAhgn
FYcTcn/s+6W/zucWbrRxkLNOJUqR8vAjQiVNXEEegnV52O1qdi13AgqLiXlajXTE
1VRY4KSHfNjnlHsye55fUlBUpUvMAeVV/ogy4YjmTVWN/PlFqOrAjN2KJBNDbtUl
bSLCp1Y88u7M9OoDOTQzkeqEXAP3EghvEyxAT53AsmqKX7mEUlvqGrLlAP6UVT9T
QXEATcnbqBCq7CvHa/1u/5YZUj2mPEjyuFPAekQSth87kikAJsWOqxbbXogPHCau
FJFM9zRlleRGKLs8NEKjeeiLRvq0SHQvDCuoW+LtHmFJpFmn7bMWD2uykMFbY7Kp
moGLLk6yoMzKjolHvoIf8aNan6oFVlYdk0pJOXuZ7uWd9S/cPQiK1/i8E9u4vdZ6
GIv/2l87qmCePNt3h/K1nMC+e1LnlN/2LxfzpjTQ4pFVTpq5f3g7VoeOpP0w5jDn
lxaWfVqa9sWZ4WS2hhO1BrdETR3fXyOMbzt5FyyhBeB3jb6pzvmttNNdpJm8o+j2
y99/kXFM2NdYW3uK4n3VAGF/cJrjVRZbQzy07ghAtSRxPqMlwah8AxzgnrP42pUX
IxrmfpWgenCCtoaM4Y6ZztgBwGo2enz99lJRetaw0EJiNt+O0ZfzI2kRQBHEcdzR
ydQKSDvNBjYhU+D+4//4qhYSFfD4cdJMhR5xiSKAnC/+Gj2cIgZpeAAnfs2rUZFT
+ZUJHhKx+iBeJVCEPIXv85g2qzn5D6tlWiiSGXejPxbxsyJGwQaVi1wTGfZHSzTu
84HYgmv7fVlKGU01XsaSiCwoK5UxpNC8GH07HSj6EEYG+l8JwCGBjAmvWVuRdmgi
Yiw57oinYQfx2Sg5lEWMj5iilNoezdg8GggEDxSZcahtxHBf9hWB0+OJA/bDHB2I
jEubddqbpuFLcpw1Th76RZS/VSuWLsXBNJOn1IM4u1YAt4h1aCG00Nz61XuQaqRj
rsPtTDkwjyO3U04d/A8nnZXqEAxzzTyesfqSaZ+o8khtojDPY2GT6758MJw5GzEz
wnmaCrnDATx2lYfSOXGjn40NjQzZNGGUSSjkSJqIbydrn3K4QTVb8oRY1dSVqYH7
4TU9adgVkKXWoUVPbshycck99yke4UflSHxqqJhoNCmmGvh/gk9ZjGwPRTNItMWc
/81S6EZG6hA5ID9O+AOb3wK2JlcqRv2BGqwe7lFWM6iS6ShxXIHPo2B8Hz0El3lW
PQcO7Ar7f9Ig0p4m+ZywRxQ/RTxOsHVhAPy80esit4M8RrmMu2GLtqOBEZe5J8R5
14HF/v74keOZd/Xzc5Pz66MnXXtKbVazFHYL6YFpSUHiXDDP7jqucd1rZ5MeM57v
S11hA4yqcK3TSLZIrbJ+slisfhtO9BHNI/ZmkEJEQxpSaHVGwBAWRnvQki1u35U3
2pQ/cW1Wed/8k17YFRhTihd/YjNDKIGOHlNHRsFg1/pJlh1d5eCMOooS0QD3/j1v
e1J/+9Y5yaypEDVA6eSIJtOp7it3g0cEI7UtDyJ2Lhw=
`pragma protect end_protected
