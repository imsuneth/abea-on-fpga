// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:44 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I2CgGC0olwMJ3PetR32eV8HoV11JDqxPCpolQ9ZN2IAjpF/vtW2j81DnoH7iG5cE
WtNMd/q9szDeSY5dggyZbM0BEy2zb0tpizNS3uRZmX7oEC+NDsMwB+hqGbtOMJGE
HxxAWOnxp4mRkg47WwCKIXS8qJHhZOmzr2DemZSvEsw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8336)
EuspwgLT+Bebkw3Nmr6BA2YToghwxcnbmCsw6uSiIHjxpeqSXGj9r9BNDWsZx0CZ
w1yrCtxcamxg+zxXbxqBJGohtO+HHWkR+ax9gS1wgPao5TOWIZJ2KwvkB20TqKpN
95TJZydrrp/hN0TDAsJPrGw4Qyp4wdEqqeMaUad/ViPN3aDv8xxsUU7fb/Lr1o+b
EgTAfwONPGaqjXLWOiztHsxTrBXWitlPS8a5vf/N0SwzTx179iU33HiCjebSKuZf
rXoRlyeoiF5CBK8Ubuib1CJFiDTfBPW3MqX7t1AQ3rDpdnvQeqftFrnSAzkAsMDP
wvCpcxp4BeVMOGtfe63YGQCO3571i2C89TlBFyAVJB4V37z64skrreE9aLAobVmZ
PZMwUP2UlA/jK33uGgbjBeOFd5HkFIXjsD/NLRgE7n9nST6qaR0Aa5fNuMNW7f3g
QvZEePrZCUDLRZVrYPWaq7KmwiK5HMuHkSW3sizpf8230nwlU2XCFEk8H42mmP4i
ImHafg/3fokFhk331Ydj0jBgdhzDhLMfCzzdzv1A1Cly6nTdJCzn7481gn9Er1is
syGOlRV2UsSbLvrAxLAlEn+tKEs98yFTMNUxaDHpR1K/F+QgRkaIkaNvhku25aCu
xtoqsLT0QvlcuN/wukYDlcYXL62kSpmumFfhyITLnaZTEICQ+aOVZ5c2v2QIOFz/
YRn0aiadCczMM4Tz3lT86LvfvD5PuQME0zfmYYYbqqDy62rR2YmjHBrUmfmwZipc
5NdNCNHMIaPJDyd+Kz9f7TqFRGDF+dV0Xg07I9ziicU+1Nx3Th0c+/MUwg9uOJrr
YEGrtmnhnq8QrkeI0g6y/GmMM+rQAcMMf6Y03mddcU1ly+VZFTAzB6Qe+mgLpJeq
Vn6HJcp9pd7epga1+ep2ptj2G5++dSwXAFzAPMthlUXKrdC/8emTwdDtU1vkx7v/
ehebov/YtJ/SRGhPOqDX4JF8Lh/KQnx787VHxnZ+R0pUrMPn4WLuDD+j2Qicuplk
ljoPGy401Od7gWRV6sBxhLMbxVMq64G6AmgzMqzPX83f9kpPaJ5QYV4rNPAUM1Il
c/A2v5HTMD/Ta15YJQ6dUe8AyBgJpQ3lRnASBEowxy5mchhnXuR5gUyDgtmLeQCs
J/Zyfbr7adzFuSD/TU0oR6mUbktJHBY9BL63pqf7gTIEzoNIKJx591KQLSsTjaEt
W/zt/jef0YHeIu+HRGmBSTwRjigYw/+ymOHpo/8hp7hKO/g6s4a88+eDn2mJ9X/n
C1CBxVHn/dNQyydWJgCchxirehzDpY+ziFrQX/t+q6FTC/aguo4zTo23443XEkdj
Q2LlITlKr81Nb+0IVcKlvv9qm+Xdsqd3FTzcFIOfZPRa6+V2na/o5rgKu3KrS3BT
s8zjWnpEgAw5zS6XUURJmWrWADz1ojSYS8vCLh8cwLak7xdT/pFnuqEw47ClDN6T
ODivRxlWx2iFly3qlEbmqsECdZstjpzcANXYX0E1poNCZ9f67dosp8XkqxPtYZij
HHXlnyI5Ekdj+dxWYtpBYupboHphQ2ZrVC712qHOxB4JQk0iIerus46UuUNKmV4R
sTtexA45u7/TJC4pJDNmmGjY1QrVA59a6eufDE0d/pOX8Nk+VvMBHeX8Tv6CjN47
zKQG89JuUIsAREXxtxwwA6gKaENMJmJI6yQdHaYoJ8qpHlqHsTTb63KThyAOdNnR
DB5UwH5j1IRLgN/2U7qs6QDvxMvIL0An0oDUbGvn5CcxKcUhaeRxYsQQ5wXqaK/q
4xBZi+slNyCToASGsxopSIT2z04aSsFBAi+u78wHVA3GxbbBQkm+426k0E65Hp5T
L2Q2+hENG2FQCoc3Hn5GdHdPPB9eq6vdhLEsuyrFayHQKVLJWAecloIa8QjqSoGX
aUYHmKkUtMDfYqj6rlAbwqBaJf4Od7hhAMZnz5WD/hhrPujMXknnGKWJM5G/Ldik
N/s7sNDl88FCY7ByqKuJ00T8s9utf5v08jI0dOFqgpPEa/483ZCkzSu+Z9pRp+Nu
I50aI0fEegXZ/AqLuY1b/T+bEefHZJJvnq0/8sFmXNlXg/0/H9qSYthVhVMxS8TX
/IIqkZbOB0pDZqY/5rCmonqMQ9iGBwncyBhwzMhFLOuezjJqimvg+4n0bDpA9iZy
Ow4Xf65mML/9QyWrMRuZMQFgVUtx5uOY1R+k2ODI4C/+BacdmVy9FC/LhLBjpbmy
JcMz2DQ1ctBh0EgafLFCTOWODJHmdNIDR85l2Gx/FXFNrxsuBi3K5uSKhsjQI/Yy
5I13uedSMT/X0bA4NaIuO7MDRcaxpJkcTbwzqLOp7vlM6TIfAJkMkbViG4Kd3pk7
nyT6gGTc71gaooeQXx00VxHw+OQJqctUd/b+EjytiZnG+ENTO0HgTkfJBkcLqQKC
D/nPUN7sum4wpvKspXDymzMxhz71iZ7Ln2g3t28H/njRB0ioL4G0wPBvwbG85PJj
VwqYrxzLm8CogWuQuykF3ustN0LRopnXQ6y8ZRWA0S/WbVkusUTrh2QzWvBE2ezp
LNDGn8fDifcYkUf4ORvb6KjgZ2heFM6iINOG6jbj8k+Aq8Ew+62GcTziydfCukCH
eTFSO1MHuXGHQCwWin6udwoTrILyoZW5j/tkDl9yNrYAEfTFgXV5G+PIrSDne4hx
gQx9riCbn4AGIpRsVtome1PNc9eH3+uZwKcLqLcf/9D4yUTOxCxW0M1+JNZoj8/g
gfd62xz88Elg++00D54J0dzk+CopxKFGioxGpA++Gi68Y4NlHmCfWqNH9HYiNncz
FbaKYf/skxPGKf3fBiF2fZY3mWL9GbL2k+gmd3/guJyBeoCv/tljw90KN6Q/4XIA
jwaag3oNt1gXpMjF3WTnel7+bR2iBg2776aRg1PJBLlS1qko8FYym3oLckRqR5yz
1D7yUC2g/LvF22wr7NjKNAFGwImoSLOkAtg7JxpHw3BsiUlCGnal3KthAVl/xlfq
kddDpULK50n/ylEQTgXJQUjgJCGUv4EqScv/TostqeV+V+eTCuGwWWXEEtULYvF1
y26i72ct4xuBOfws9oqVfs/oX+tEoEL2hWtTaCTHDV4EEnBSRFxijVzeadtBi1cV
V+52QTZlincEmaR5pwyt23eAmdxiWZz614tbKx2p/PCQNRPVSDMoYmTvgwApaw+E
cTyzSFFJCksMvnILhUOy6KtECjxiACzZRx7U60A7X69Q7Vtn3qsk+fSpf4C9uiX6
Nn5lNpdx7PM3ZPlRwbxg+5ubtQ01E6XJR+n/izHlrqXRZ00GjjuNFjsoGcZ3K7ZD
nsWavrYUXCVMlC/MfG6jrrM1Qi6BaXFUKzxg4xGPpHvH9/E6IAhZsBYe57+E3x4S
ui+6xDEXv+gePYSkuOxX/TvYcI1Ri1NpfzASPDpGybflQ7hnW5jDaJnBeqf/Tohb
qnI3v7D4lJTc6qDrWEqkbkhm4QHsoPdz7oj+f679DM56VvoWQfpi+IZcQBgA5bA2
q0rHdd/M49qexvblWZMatXanMYCciGRDpOskIMX8ObESaT+y42DhSVJRmQJMA05d
G+PDVhpjsbrfmiD9Tmpj8SxLUsfaSbVV8arp/lRrcsO6+18esI+HYRllyw/s9Jlb
L7kOJCBJnyxuLOf6VlxAj2AbwZGoW5RESUdtNymSqfKP0wuFr9/4/AMnzjfRhb55
qq/fvbqgoFpl1QOLUGVL4DB/YKG3wUnKkV+Y1eoMqLWC54C5yevp/xYzt6wizGJV
Nyd/LoPIUB1R+wnFS3WMcD7cTn8W/eNDNnB5QAqO0wSnb/L2nBxQOTjMHtnPK5qi
ShX761medtF4BV3O7rqxVezGZTX4wj/7mX6Bbydn6KH3H/uAewaGmVmKN0i5Nfhk
9V/yqu0LK1SD6LaguR7+C+920EvFlt4XrZpP55L6RG1RcEBxOxqp/FZoTp3x4ZxR
/ZmzoITCXQ3q/eq0rjAj9d9Rfn2xNMlFCWqdEU0S0VFq5+AP4m3+/TW7GYW7wCzI
cZS4w0A0doxIQpt9Dz+IShJBaEq2KRP4g31f9px64LpORS4oycDRe0tbXok/5O56
0T8PrKwOyYUEArZmzqEFRo8YcH9IzkWsIDDnnxvAAgKCc3wc64b/I/V+al0693it
NlNzbIdggXFB7qL3UpRtLJAeIpye6Wac+Wtq02k8F1ZrWtY16Jgg/W6976/9Lvqi
T2Eyoo4fIW7eLvFPMXSbX7P5uUTAB/3vvfcTWxnGIvXkyy6+/iCBNEWZTlSTlQDa
OT8iYWq/nwiaooSIMIz3+EMuX4rl6Bd6zTw6men2I1jsl2pZwTXixN7wMtiFZyev
39RIjt738zP9rvY0IQkJoQbvdGoeHPn/fs32+Mf8A+UB9RN5xHjvk8It0r0YdBov
VuEoDNUEh7N4FVm4Sp6WRpJC1TaSKqOKwy17haCI+bbUyu87pHyWARPRv2loem7u
ER1vX+rIhjX/wZXsQxhkhzVxeb10rbs3GUeb9n/au57m7LJqdREVbAUhMwOElHK9
iSW+qRsiQgfpAhpcGbzN8obYr6RcyIHnNlFt0xk20x5C66NRUhjeesosCcKyAXZM
i/sKdFyhFdxxv5AqU96SJZFeZm07yQ87BQNr3FSkM3iJ66i7yIld8it5ZOYnOKH5
Jz7dYiEeI7PbBC41MwCy34nX0ei65b8vzqeloVoJYbrD4O6awLbKr51kECAIawD4
wfi4vumqSRdfH6Zjz9T1Z4NuDVG9yhv6MTT/nU6iuCJs+wM6oWCVLLShC/lv5ln+
3GgogCw5Han3TcstLNKpvetCkkP3Qfvb1qHWqrpqdX0QpNrSA5GC9FyuU+194Mkw
6Ob8BRil/WDCs9GszytUmR0M8qUpXjQN9iQMMCgQ9Woo4Bypemrf0EykgSS5wyGt
3T/wAmJYmEAC6zAKWwDGa3XQ75sIhHfZ99PLPU9Vl5jbsafQkXhnJZemWT6Ajs3F
40EBb/NUu0FGiQ/5bAA3Md/cZtVEGR2hUxoaqE8e1aXBWQauA9+w9mN78z2p2dFg
55TBIxOSCwPDnZ5ShdjosEUGBp8fJR6tNLrER9nRtPqnn60X37Qs7FH8ix14nWuN
yyN8dxyU+NObtq0oa2tryOUTG12wwhuCIU1tI/FKDxnbIH5w6RUtO0uLHxRy6IYk
/nkJZE2yn4xjLg3r2N4Vg3b7pss0cKlYbJqpi796HENeyrAhjHRKEy1VsIgaK1Dl
6+lLd+fGPQQ2TBHVdFWBTjqqIFevxqOaXxhtBr49zeqqK/WxRtTsm/Kn4syEx+jC
2cr6m2C6yQw26joVEFJGp60TK4Ho/Pta+02K2+yN8360duGXqUZLsap1oDTvUlv1
Eu2D2rOlsw/iecdlIEkwlRC9YeoLPVyQ4A1RiZXTjryg51gV+Dre/sv3e1wmsCDx
f466h+b8EkwxnsQhFmBWP6n5g5PT83cvSOggKTs8nKto0FWMeZBVjBNca53BJWE4
1S5PWsr69oRDjmLLQvftYi47i3CXA1G1zKHmfFtyJfsSurrYv790U4BDVjMYO+dv
UaARmmlBqYbXpljzyxdboA6Hd6zcJG2LJwFFBEM4UyfcnNiAUSGaVi+lioxAU6tM
xaFu9xNPNVDWZfPEBzLER3V254TTP44L1TPAsCa+1gfjlVJHB8F/JmLx0aslUzb0
8JQn0+JD38brweSI8+qJAVNxv6EtU2UEm+cdsQBVn8YMiS1KfiWGVd9jdZyeKTcg
9gh7+CFmZCEpPFFEzSAIKT36BoK7JyhdxucnlAOtkQWzhGfzNNCCuLdP2oVcc4i4
4q/bGnex9CeSsRSAS3HuyppGYxwWhZTbrOSrIu/vNS33H1LhU5ALDzMRLAUZjVt2
YBqb17Np9lkTsbx6XXVGozqLawOLWaxnazPvsHuCQBgNn87fUE6pRpFboWlCcHAI
GQ//f345PdKuMmz1KwZIplF8rq96ufxSPGzB9lzK+AUuFYXKL6B5bpeDfpu0/Czq
peEVdsOaDeWCdpfcazITyKk7An8ROPbPY5BVjB4F/A7F6CjPYzo0lUss2X3F1n1B
wO5N4Dr/h8iYRtMUItkirx24npZWxT0kA7mPpS/iRDffytvC/AfgcH4rFuk7N1PV
5mh7i48c4GG3GfyqRDz3nFfMlNedhclY5tE4L0jt22FrGk3ESUnPuBInM0SdpL4y
xUsBu4kgelOzLLFRJ937TYO+yJyW6GoLV97Ar6fHXGBLYUD/8QLF09eobCj9v/U2
GqrNqUGmKFvmsEmzJN2we+puBFwRo1qef2dZx/ihQwjBOJmum6ACtSr3lll0fbWN
NAxMgtShQYAAS6Og8HmyH+iz+Z0R8IRxmPps8RCLnmcjASjXzXc47Qj8U59a3d9L
ojB+NSoRV6Sf0QjK6TyDLg/tSoffbI7r9PMXyJxm0tBtSze7lfmSmpqjQXAocBzC
xgviH4+jMR8J1UlC/MwZA/eyFBarPaWPGS/hOxpoBUfAAZKZkQtSJbQCy+0wEcKq
5yVK0Mu7RGyCzxtsSkzcwVJWdwqg9mmzxekPYAVGjhI8Ycxo2eAdumJ6zt7ydX29
5CKMisjsCl2h/fKCQXmKXsR0uKXz5PHcT2LaU3NtgLtAiG6z46NLwIIKeey/JH9c
TzD4fzN30wLfMrmF/3/PyeySgza2NpFFm0tPTwAMNLj/uK9l1Y33LsmXnDQ4ThkX
to4KTdua6/MfgigUhlPQkByHN0jJJluZpO//cPFPNj5GLi3a8vVahmHTZRR1CGMX
qAx925By6lBkonzXgN7QChOR8modUw8vYZ28ssDNE8LCGXizgeadJ1IloV+nI2Aq
CVEN1ZmNkAHu6/UjwPgbHRYGmMNwOMVCG3vtVteU+2k42LxHLJbw6JIx65sUvaS+
evZvU2oW0KCJg0idkKKxlChIkaDI6GcAn8h0YCwNBlbMJdsW6yCQtKGBjxwLQCXk
+TFm7d/m1YMJfp01GTWwKowoCEPypAhdmjHA41LIesrwSIUw1WNtzrNdW8RKJKhb
vYpxHAYMoLU1/GAPX9gYu3LQF1DzNA2N5Vx7lMlSh2BvWj2OcMORDPSYuNFtQxsJ
4e4muFhqrRM0gJXpbOftENgDsKgeO6QIusRMf0jwJ7vxKKRPnumhCmV2jiwMAh0y
s+xpVQsu4Zufo/w12evAwFZnFFpvbiRzF86XfdQOZndjZpECXybw6xy8hThL0gWk
/LOBhhCPxIa8X8RNFfaRgTFA2ADVaKT1cKU64+iWYVAx5PeuPmIJjxY7dSgdCABi
Xam+Xq9gkbzWwxIHClwz3RKguqNFJfhKvAEOPwjSe2UdFFxoeHy/sNQZXHymp40g
dE1I5DPSCKqy62oGqHf0AiWllpGshQ+4OkJZpSOXv96oHI5MsUulbW7UqPtBrZNi
9w7buTvl+CXkHgWs9jI6qT+5kfxIcl0jH0x2Op4sCAvobPihEIqDyurKZYpagLe/
HeGOkCm9S58o+fzNa/+xgi3bdCvREIY2E2dD7lhca9f9rJrgswfTDfcEkdH1Ehnr
Y34oDVhND9OLwbmpAzUR8b3aQDUB0zztPsxU3P6SzRKfd/u9PS3Otpb9nZuNoOZS
FelXoO9i8BvZM4q7fz2q8raLMi5335xDMJ6yD/eShquDK9avPMEtJ0Y1i7ZRhna+
KqhRSP+rQDeUebrW0UTnEG8SZ2xjEwTrt+TcteYie5a4hs0hywkkpSmDclOs6/HN
YgTLe7D1c9spqUlOb4mSLNde8qrl25XkkrGoSJmClSgm6qQkxUJ87rDhSNYkAiEw
8FgYm4oBK5aqvuUjANVYxCF533mT6kRh7Tvo1cjWrgPxTRGzMnETojcalCSHtrzp
r1CssKdBq+HkkJSmny+1jO62gWB8V8IynbDnYTvAz8/+C3k5o8/WaF7kLuyRxY4R
iYPL692gAkRUbGhG8d/+hCgtCIc5FczHMHSZNei0uXMnZE6C73ev2YjK6JNQ4PPL
DX3sECdETZ7W/43KUjrZ1oomYFgelG0/IPAyDBpiX3FWcUQ9VLIZDpCpOvRgNpPs
WM5vnz4GXgFjsAZf9oRP7z35rqAtouGmMrKjB+hfnM1zYhuYTviKKyzM+wvhvNi2
mRdcYkz0gvr57SykUJDQKhudLL2HxAwdmO68dOs1rLgZ6HcL2P2tyZOVG2OfsBg4
5570DrDg7SkSQwBGHvS65L+XjbPoE2lCMUx4G75HEFERmPEBC9/8FnnvHxAxzCOV
XcmqBdPI9E+bUTkHWeok5gYnHOhfLcdcAmRRLB9Xm2WtjYSbisuxa+BDQRPMbWCc
2bBgb7gnHdCUYTgmFlE3akn6em6zhY1QNq6BDyK812Cl6CV0Hf38fUSDTLDJb+I2
NZGEVxsOJdYRkDu1fFIKBnH+qfEmDzJIo4FpXIby/q6Kxr/pwC0LA5RFSk+ZgSIK
ZZh5n+3aSUx8PXXwQJIr5IUbpH+KcOLSlG4PvQ29uWlVMGeUCE8anhMuSeHM7Kh5
u6FZBJmwAJ8Jt2R5RiAy0oGhabfRpbBaJFpr3+TiRc0+QeofPk6hZznjOFpb9HD4
GwlTaS0JyurButPdBw/wK6N9f/t532mPIN31SIytqABgh/pdbWE7dnjEFEODfEU3
sYZPvYLWvR8fJH3WW8/c2sdaoLQB/T/d/SfTdl+tm3vYQnIGYSFarHLZUMNvfQPD
R/h3rgF4HsxHqzhhC2yMGq4Iokhwdq4m4cLHSxzmEXVuCi8SjVYckXwy377h78ZP
bZGz0BaLPPSGqODot5aT7ZpyfA/mHbfOE5dax7ISCYcKzRUpEvwEyIDq7TViDfFz
AkCcvAKdhrLfKl38pbLjXhUFJ1c/jKpLX5qGbUxgdEhtkQuL52ui6igvKofy4Saa
ZcNlwv5Xk8Fz6kkGh3CihNgTzecqrDAomQOehqIX9eVl9cnv2BnJLyE3+qMzUrYn
Re7n9gqqB6rNAmvvmD7fA6Bk7yI+NAm1QYogW/d56JbKbjJRYy2HDAcLfPDiNXDo
gtViBR9jFpi5NDDouistkv3CFvrtpyPbU6N1fa3rHw5SHOb1XmMscUS/rUsSkUNr
cF+inb3Fs1bfntWyTkoa/nO4dFw394jbWm3Ep60D0bHBhKFEla+BPpmmQAAthQ2S
hz9WfjzObwtgxb82Tew/lVC9J+n61cDQ3z8YSVKFY9A1omWsTJNcoubTdBRiyz7e
aZYwAU75po8ssAOyaTDkZeQLkspJSq82WQKv58qFbFGPMT+TSGgR/5FKP7ZG207X
33T6RWR6W/i2zOcQCWPCGWDFo60xAcww0tY5KE0mDMvvxIRsA0/pL0CplnDN6uMI
KE6LgfPZmZJqZQNR9H/ps6Onz+CGbayoORpRw66FzaivQuhjrFQTS9GYmULCKx3r
V7DCLnYwr/WIV4Tyi30eNDk83O+z5amW1tTWfa9dUQrsp0iMPOcJ8tFdQEARLv73
aPKzNFOJA3YPq0OKbZscFUcpF75neEFG164yzfpr3fx0hSpqf0gSoMJKqdRaPRuy
6cIlXTLXa/wUGjlASkzCYC3tHDINssRQaVFIl8DT4VTyMMj/8Ad0x/5Dl9abzv+A
8XRQ0DrGmYuXmiO66my+/GLBNb3Bbbc9aRjjNua91Ekj9iEEo5gAZt7Npjeho0Pe
ClyjgA0DzlZDKHfvHI0Sjc9HiwFkClcBASFYsOBVIOqF7tx5LWTiladvvTclZCwr
+4JLOkVHRRcrH1t/EztI0cGfN6noKrEbfPOYtIpMPQJPa6xpCBymKpIYCLaWUivV
mRo/tJ2Bw3ILyd6l0SUl6ONR0zgEP7XYV3KhIuOXlCur1g/DLkNkU3vHFtK4G7ay
+3JcSjmPzWIrzjxgymOn4zZm9u6RMBIDHxsxl8pXL3Bg7xFRNiZryGrwYx9kTRdx
rolqOqOPJGnc7ZdeukUUx+vvSxs5xkrTdRm6EBsZZYhij6tMA1Batm5EMCtK3sZK
FyigdA7YsAeYwZ2Urn33lcl1irvQLCjv5xoTqLRlikCrHBiaT2KXEJB+wTejSiBz
cQ+De4hNiwNODAyKvoUroxKNExrydslmZVoJrVWbQBTk+gKf8fBozmgnoTwrC7Th
eGDD1EKQaIivBoExjk8YHmec6yGhbvVBqUtaXEn9HPsmjxFAUEVmjlC1iVkOW1jK
t+yzDgVhpydW1L8UTa7aU8bPTeCWrr3Lbg10wm9Wo2QhRL9Xc6IpQ1FD63Pm4LkX
u8LrK/EaPOFqnz4GbapQGWO5zBDzv4ehPmGh+sE8hbZd+Qjbez2q1E0OI2LmG8Zn
EHM1bYXGeXiVd7kYA54xc3nq1TWGm36xIp7/LJJgsw/YXy4qQxswebaiskLZ6N4i
02kgI1ioG8ceIsXwWVVJv6Cyu4Hb9mbeOcq14kHRYuPy7FRKJq9LTaY9k4cQnub8
UsheE+H2JOKcTWjE29QohpZRtA4QF5WSCALm8d3/0Ct9njEYt5PKu8VYDb93rG0N
z3NwmZi1cZrbKXueeLXfzbvdrDVybDV2PJGHqydJ2ReT/BMVynoKj9WIT3MI73ah
/KzihXGE9qIyT+aFGdGYRFOy8AunRiUUBcSFTzyWpRpO3ryx74jXi9ukxGEBY9Fc
JjTDS9OXStZ70FS2TSqUi9IYM/0OM/SFq4Ot+OCdjXmxSqnrhz5/+WtuZ5IUqfms
+dfyghgyt+4uWRPBo9YmjN23GQcTdEq2t/N1Farrw4naoqgXXCVNeSdNY25yCbYu
n0cxBKKRLIXFSsHt7Gy3pN92CaIVlOMVnjm4wwa5RuQkmAZcnxt/8HMx86MXIk8P
mjWlZ5aISUvGKXbndC7uyncbaHbz08ieIa2eDGcxW8VTiyH7Cmtzzgck1voCM02U
bWJfVxxcHXBON3q7LTnDMgEhahL/NJzTTfdp/AGnwv3S7qQ5dZmPa/htF0FkftsJ
V4c5aSgRCXSPlvqTJ248aD7GOFH4KuBhMmbaMMRBL9D6A9QWYs/bLBFN+Q+gw5Ht
6fseZDn1saei3wQvpEJzZv5q3HCLtZIo3dOwWAuCZgyP9tyNbthzKIscrdXfjO+/
E5aWEhQDazIOCbAhIC65FbylrvpX+39uez6gcyIla7U=
`pragma protect end_protected
