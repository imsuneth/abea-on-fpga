// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:58 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g7feIc/JjOTjhHsnaIFrB9gICca1bCGXlUiVPdGedhAgfzqlX12AascpwV3wxY4H
AQl1yfNd85SLqy0KHQfOaqxm3bb9hlV+QbQ43wQPgp0DU9lGg0Wl7rZGNWA7VoZs
LUBkGE1md/iM8VC7CA+a7qQeXaVEtGGRGjgmhIMJ4kg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25872)
DM/qKMCvzeyxIB+jRflRKEf7BNouqHHce+hpYcIgrVjSuueQqTNMyeQLo0twnjvc
vO52kl1KiOvRy21LCO1rAA0lJisO52j1co/nKCgdov6hIme2qMWh13y33yA5+EmT
FDcsY+7KrETGL6ghhxrCD26ZJ6yK64oYpIoq4hGK6ecQ4qexPz2wdsx4r6wxqZIE
Nuw54QXIfgCZRBUmF1dFtvt88QCV7o2ikoh+YtsYLx7MdiQ8Bu/HSeJd5LYIvNVs
EmI27VjxIGI2ds96EKir8gl/rbJstXHEJMuwMKaFDZyCgusD/m6QYyovB3IuDbsB
tZbOrX9djv85PzcGnjz5tUHPxgmAIykmdM2kNPiNp7DgIiVmP8WuzwNY/rEEPsxr
FU9UWwAHcNWjrSTFeBnm7xDF5NJUcd3VPMHS77o9yDKDX7XbGrk1IKiEFhrPhMGh
rL9i6YXDJg9dLIjHRPXOdcpzvAnwIHO8KLWY6BXFG6NhaFzwfJeypHAle+Gn3FkN
vRZLsaMRVe90ZZGYdoZKmWmVMH//lpUke9eZ6JV205B5XtouZZQqv2LlOrQ221rO
hdsU/8JCEm0DQzWd04PktjILXHRpcQN9M9yqIygsz4ahtPWczDJmwaQon/OvmUHq
+23ercbAtlC+Ad4ypIgx99wzE3undjGAJt+Fs/ERcBdT7KiX0FOyVb7HG1Zc0oZN
C/7DRvlYN9esr0QqPP7CASfCqY1CK8Nc19ftzUkAPssKGC/o8ze3zPBtHiDqt+LG
FDNa+mSF2lZ0uSCsjFem7sRTPFSbBtoZ+zxOxBm5oMXFnK71pPSPjVF+OamVZkKP
11QEkotVHwPaRkkrUfL1nkTyIrRQNehijK05u5oKQ0Doqza/1PAlC3p8ahs/OQU3
3Pxp018pPRPlkDHWU+rhPYA4gWd1ZpfuqlSCjy/tFXZ5IYqrYtQhEB8wpSZZpass
yRrUW5TOmVYPJMKZJrE4kme3kTiz/SG7rUHBNnxZAnvGgPKlMsbjn+T2XyCefrSJ
Da7KevSNcNX+Bo84Y7Dl4r7cBmqZKuBN9OCE4Uat2Fz/xLtiIQu9aN5/L84W3Vbj
7BBmcGiE52blGwdEwfLmyqpr+Xaj1D0Cn20gGDtvfPMfFZKIXeEH/r3a0cAKKNM/
6qrevZZ6UQjqUG9l9RnV5Hwcf6vcRsswbMuRcWgP3OmXVN46PsQvVLthN3AcckFh
4eMCEXi/o/C5A6amCLCsClIKM+RFHPa3WNWxIoMuxyUtvowN/QZBoElrrjmdO3Mo
dVxOX0qw2lCxb0P3NrNQTU8suAWPFbZhqolOfd5s7Xkmw99g/TmfQcckCqBiqeua
RV0IdhUsuK8XLqRRkj1syHSI6ACoNjJx9erSLHXriwCIP5Ip0IZr2vDXK1U4Q3Q9
HrpdeamvD06Ny9xhoScPxSKnAFOX7GGTwJN08dAn50l+znd8kmUJ5PKNZ/T4R5+2
BacJb7+uNKt9rz7X0nZ6RR50sXCR8Lfjxl68VTHwjeAdV+i+Ciiri+c8sAwsBx92
+0GjgerDJlYS/aZrm9GVGcWHlA4ZeuRnCGbc1nUdPQVqF5dPvsdRDUQRKcKM8sJz
XZ3VU/2FJ9DFy15hP63OBCZO6Fut2O5nyVq9WS16Cpf6OX8NnW9HId1UNtdjIbDo
0iFZXg32PmgL+Tg58tnyw/CSluExOwOryD9gpmcV4vj8WUu6CHpv0jM3fOeE3pFg
ElYfk/31sPEiq19AE0fTdMeDCd1/OK+FvrMSIY1R26mGDog5zBGJXM8cY093Hudy
4Dt8oAL1bEXdH7ihh1QSM/ibiGMJmT7PLWdwWTaWNuGfUaKEQDx6fU06UFtisJQH
7Lrsv+ULxG62P6GzYArgZIHEaJYd7LloX5PGbpf44nKASrgK9oHmbGp5d3xXPwyt
LNSAvpuoZs8CXo1Sk+gwK62URaGtC2Dz44dwLElkrJ+UwBm4naK3SUgAiMRpiiJq
F3rC9nHNFc1XQ21yaEsrF+73cHd5Dp698x5MGDH/mlKSiKJYGYMZLJ1Ee1HmCTRO
9/rkjde8oc+hKt2XqlDC6He80SQBOem3txJOeFl3LYFPeF+oi097Muyw6mfOI36m
SlIpFl1a8JXZhbeWhMPx4hVfwLnISu3wKBrf5tztvGUx5Wf7DiF3iyoBzEPDuHtk
lHQJLoEncDOvE7uQjRI3+xkMn3Hr4MzycuFagsNB8mC4MvJDO8naHJyJfCMNluns
iyQbPPnWQxE/2odnkIwPZfEAhuGFjtymQuFJj3SoIdfeu1vCVuWALMSLcSbvcwcc
FgDvCH0kxue98aUeGx5Du0gCR5/k6MHqEz6F0+Hcn2kdYv7OQknI4Ws1/cCO+u/B
uckeDx5dUlXd+mtminbgfA3F9v3NXZiXS2Ts2mN8/zB3qcbX8L4rweqKJ3foWfbK
yE2t3JLsVwpTOZVWEpzy8Dv8Z5Ug+hN3vdu+0oADBb0HVA3wrtTJZgHmeWURvHtf
lVgiIcqaS4D/FbspQsDaej+AAvWF2sh7Da9hpknM+9uioGBDQawkQ30iKy9HtNJV
LBNhPG/UOomYxK3n0aMaQZwtCFsAUk0CGU+Ofmwe4AG2NTKPXry/Pi7mR3cb4qv8
bW94nHtWYKfFw+CquXIMEeEtGsmrUbRy09LF+hmvZk00aDGVQDD6zbHvjefqTDQr
jXUashRU67R43vos08V1LvmNSxp9YOydvvFwgiUcnM7ZmpbkoeuSe2c5HbewiLHT
P3dQ1mfidBbvLG0Gv0J8c92ofgjFrecUBxftTioes8R8iykXTc6PeUT9jWjFa58A
QhRdSXu6Wx2ytgqCa4dRnBotWKc8zRImxjKYdUL+pxu29AAL6GdKyqhAHgKpqFKU
RMqlTWA9/zVQnFO3JaDae+CY9ORuQl+fOTKCqgZwoBETCPPdwCGdV94fgKDBguL5
ls4f1TLv9mCgomOl74QIJJowH+rwbgc2UZ1OFjbNq2DFZxcqxGZFXxLaFSUkmXR/
XqcgY8WnDmI0rpI4DG/uQti025r5ZrTREm9ic4QeIA82MFAovGqFDz7drH1oKpsK
sUbzaToCgZ22f0AWnaj5A/gOga08wPIOOBqqktqFWT5FnokqNYlxy9MoWSdrYANr
rwHJjrilv0afWX2uypFVljg4HpCBm4+6hOeOF+j3cIWfTEY87+unRhlOsKg0dvzp
cna+r/S3jYcctKgR4fbIdD8Aeo4KrzyZKV8wQzOIsRtwgyifoEkfIfP+HYXKW+WW
1FSxKebMpvLMZ0lFNYGwEwj1UopJ3MVWaDoK9Sb/lwfM7QN8HsaXxL3Dsh14mQGm
fST+VSeFpjtOE5M+eXrnuAw3d4uBy4UR569W1B8nAXXnRmVAWUkDmSDtuAPRfsjT
8fBYahymoC0UD1sIGybY33AaoZZcQufJ050Q2+NGgPBuWBzxq4dYPpCPqrgBaFIs
CdKisdTKD7hjzq01kPeBVvg8JlEG+wTwHTK7tae+uielhlnUsqK6Zsj1zEZ4xmP+
p50xqr+lEIEmbgc5M/4sXHQHKhMZ4BajN2GDishQ76IKadskGmKFb6sI9pM91Gss
46+gZ/hVnNEWzZ1k99Z4PxNgGEAkKXcahj+G9YYpmBtS4JpYCLnke53Li3ziJ8Lc
PAeOjPN6U83KT2BsbT+Rpv36f5LOtyyezK9+8Tvazbgke9NqcfBzDcR2ltn3kGUj
VatF9oQTMpZ7nIM65EmTPvkouKTXW8HTPf+8pAlBqIwcJ+WS14b5TA4mlxn+6vzj
P+m4ogYoxY399beVLrMMJrgm2YGyLXXAPr8Ayv0PRWpqrQfQRDUv2qZxKHdT6B85
1rAoBv+gPF7JomUVJ8Yz76G4O65LcAPTRnyiQ4h9gjlXyN5p/nfrB5LNKSBEqb6P
VfNOp+cqtHg68GeYEMopk1Mtl2wFwb/D3nD9nImYqgSLYWOfph7cvlGNEXSdvmV/
8awTeIim6LU4aO3dNSbW78rXQbrK0mXR5UEMOVG/Z7FXC6lbtC8Jncpqau6cCJ0A
9uZzNEDY3RbPivZZU5y3rOVMZNmCqoEhgf57wQYxqiZGwHqDYySxhzaIOOGOAPBB
n+F9f6n0FIh9geTH+kRMiwmrAq5vGvOulMpClYIqmc1EesNEB6qJF7JBDeyG8/k+
mYvi03MbcrSpvGeaSvzKRe3sxEYAak4LVoYshFmT+gnXOt/2AlSZdv6m61ifGF22
2yxl//19nGFXBoZJhY/dOe5GRZkpNZc86sO3gdVsqaJ7qNtdtKT3XXdEDVG1NTZL
PD5nngRKBNVws1GOosdizcvzwNFvHbtHo+swUXQsQVSMf26tZ6n/IHx531RgLJeg
e52QxMWT9N9eQi3sDRdNXGDcG3bYX6eyksRO3Or8jESTQILtnW/+BUveM7EVhbGE
B2h575KS5ovBI295AQwtIalYU+BaaYYOqRsgHEU/E7TaWovO4h+K3pzv5Htb+rzF
pYo1lRb+gEttHe8SagjdqGDtoUggQoMvKqD8KLnCrKM151MMvlg8pzhYLkVGhHSA
OIRwsmWLmoiQJs0QvPewZSrcjhVuMhPjtjuByK3BbooXOq1oXEYA9CA4hNs+nuEI
TNhT4paeXd97Ea42e55CXSjuK8xJmeeoOyML8grEW/CU0PAJklSJGp4I5i0Vcn/5
VFAiHEXZ5MlvLmQtsYY/dm+7GvjsoBPqvZvWpaia5rmU4Iq9h6kdNM0QezjoiFPJ
JGcPW2uZQrmK/JVphFEcKlnhRIBip2JoFv2TqGM5Sj34V7b5l+/PG3cX8IZnN2wQ
pp+LT5CGozEm57f6sPbjwJ45D+PVcd3V7nA5yDiAuic/0dpovjzgK62V/21FL+6b
IJQOg/yGtH9elSJwy7l357qIjTeGIHSq5DkDGgICXjW+P2Ebn9SA8Slw73BKks2x
uDqN8SMVHeRCW81w5GLQSLL4WN4ubg01c9tK4qCZYOE2AzpHqI0NzH33Ovr78vF9
KHHWJoLQECAW2MXgNFUtz7gjf7zCdV9JXogPyQqAfRcvTQ0HR39fwH4R8yzjrORJ
Q1Arr+f/uBFiwqrRVvnRRXUrno1kTHpEU1p7n4VQ5gIYl2+CvkQ3kInZ4j5j+R+j
BwhpFdnZVqiqds6uT9vqxvNYsupnj0kKjy1RbCcMKoFJhNYj3tLgFZdZ323+Jbpz
8Oekvch5mMZTpKXJEnsN86DIk9dELyWZwgruMJP243LF6NQQfmqQuZb6gruDhYp0
YSWCyri/d1FRPeQtl2QXUQHH8Q3qPtZIclTsTlFriQTkgXCFlPTpU2zteysRosT8
JYzv+sfu5rQ+bV8bsDcQ/KR9kWPXJB2PB7djsMc47/PYKB4ogAMJ132BlxB/+gj0
U/K8uWjOJn1sBeq/GAt3vN+u7rEA78KFf2dOiTxMZ5kaQ1l8cUOb6E1/3MqJwdjp
SECFPN2TIlxk7x5cSHd506NlWR70CIHe4nC72w8Txt21StpIS6fPrUZRzYJ0rp8i
T/jKi2YmN4z45eNWpLxKwz6TTXDitSMqZgwdM2Cl1ePZtq3ezHgE0HbJ3gwMJaY4
E4bQ8SggsSEWBYK9E8Pbr2erwg2g9KJ0iHFpUCQ2fbWZPg7qyTZiW9UthBxW85Qz
wUZHGi8T2mpV/UV3uVQ5i1RHj/C3jFdX2kYJgxeYJYC/IcAHoWrsV+6+5vdg6Zx/
xSqcWX+RhfZr5bpCPfxNu68r2xY10tJUuCZBoWru5OvjwLkx17YX/9Iiq024qfc4
AtcmFsMCkDBqKOVZJqaS1Qra4epckMj1lkw4K5pkHY0dOraxwGIWTM9Ew8ZHOdBz
aERkMPsENZcbyqh/ONhXdTtpBu5bxy2s9u/ySsydNaJ0qZHP23TEcuyWYxH9I+jo
9Ver9OxvmoW9U2MO7tfi+DaDHR05ZOjoW0MdXxNUy9denMxQkG+DdbUCv5d3GrYl
YKfGh2www1KwT/oDcrJFNMqllLAeh23x28cWxR2+APoIM6Rk3f6IyL0uPadxbViT
xUh4NtWkRbQPfIkIR6b872a19iMy27s0JuE6eWOvbZlHa8hAgEkgELjts1HIz5Tz
Hm8GrEeHCM8KKY8xaPAgrojBKuE7jAupMi2WSpGOTW6yvIfFP41hKTrMsEBPdPSb
AvCZoPdHUSkMsjRFEa5Pto1aCqu+ShdH4V48Z+3Nh5fbVzNdYKxxY2nvmu44MotT
B/00eB4A2PjYlkuuSeBFkAlxWogBwjf/sih8qUcP8QimrGSKHFaMFqqrlPIfmLPD
q9d4bzZhZrKoOWzHNLqj/LWK4iIjaiDJcaDcBDrwKvd0FqYyxrpvYgagHIZKSwID
hDRc6XXDgBnWgzPxAO49I9mfNEuCqjtogKfdwxNj526EXxsYGkFJPPAuqOn6ar2S
WdDG25zne2rIHq8Rm5Mc8aB9ifOs5kA29u4tdLlW4iePpRSRDb1s00AitrMkqabo
FHziNU7d3PI2Ae4V+vBqax4cuY9v+aGZ3uKE1s1yGt96RMGyN8uqwDVCHV3A3bEM
FtWVdj+n655Px75zCT1f6frTo6XAnX8m1DdUAi2qqlv6mzMZ4Qfyb1jhvk379qs1
VTCVlDpzDYycs2IQAJJl6wtnZvyQ+6TvXTwGctjl3UN9R2UJN3mTuBBp8pgs1jjr
L6YLr/zaPdQTsdnrw1b5mhl6quo6BkbHE1SaN77XkYi6G5GZGI/AeUaBM2Bvqk2v
mWXD4evfhnpH1Lk8eyoBr7aIROLOfiNNitdBSG+aHdauSxAMYCCH+rCCNcffz6/W
jkavZzGQS9IV2zyuPv0EJgBZH5v3fb7bV5oiYRQqLkLUK+NLLUl1cXDSujtHJxZT
+KgigWS58b8dM2GI6quIlUqqn97z80bjEirha902XEj6D1jTJ4nAQoR2LWRKxIVW
a2rv0gf4DHpR3+9AlZOuS/37drB6u5cHKCEvr4hEGzDGqFf1NQapq4BOJfItJa7u
vJzZbPlN65rWRRJLDcnLxUV0lymyRgne8YsKFLehsHoDA93PjciuU7+lnZUDigwh
5gLTd+wRPKAEKj+wi0oLM3tAnIJRx2F0nB3Ouh201Ut/XUW2nrgcB1n3kfMR8X58
Q2Bj/9KbQMH2VHA0oA7qcvGid7Sa9+U1+3bkBySzSKq4cHzkNaXLD61TUEgXkFv4
o15KTogn35nqYOEToGYVwEpU8eNptcWDKeyo3g8drpv9zDxUokkfpykTkjaNUUYx
xEZ5RtQFnj5HiXKbdujBy0FsWRjPRxpqwEaAT4ostz3xOAZIpkekCVEZ7FGqufdu
ZB/AAjaLyJopS03rPT+EFC8ruyMLkIR2UeL39uFk7YgTM14hlxWt9rhwkxl4AlK1
9UlNhJSn3LgDFOHA8rgx0Jg/HKJvEuYdPb8qKFk8F500wmVIJlVIaaAfx5fPSenq
+/gpNnoViir4C4JY3uL11VELwjp8NNaUpIPOA60zbryyvJZKdN4ru68Vm6Jbo/BW
eijMXDjoElUX2aKBYk15IROLxIVrXe1ArBmRFnrAkEf7U3gZyHgRd2aOV9VtXDNt
8VuR/EsJnt8QymnmP/7aEWm9jRDXC8h2s0Eig8CYAmcvrujgV98CMGZJzWxi1Kep
2nhO7LuTyiTjTcookp+gtcIsMGwr+ejXuR0VPs7CW+7EFBD/q5qBZsMMDKeFcyT9
blmPAI/XCOHXl2gqtmRpLIyh+nE20sAmvQ3UKLcc1Cwm5cUJjf31D0y0z47JgOwR
bmQYySRGAJILbzSt56UbR4nhv/T9eOQCP790j4cEJRg9zH4XizWQcmowrTa91uFx
rEMugtoM/TPUJdq02rmeJPNsqo/dCcVqk37b5sov37gGkyV4H1SGkLFHlyYFv58n
xvgZH5k7pU4Tn74yfVLMnuJu3sK9Fr6NXWrl4u0ctpOfi8tcg0ksfqzokAnD0NEV
bpGEJMNJ3aqeZeUMj/3XqgpMOs8TAAtvCBd/xYVGbyFvRkZxZ5yg+QJN6ZhCRjUG
jvUk/KNPvl0O0OmkhWQqyBkypggx4ac6gmNiinR4YxhegWy0fMRa2Vlj62ufKDZe
5GrQiKlFDUTHCesWiYU37YLNSwF8mm7IW2wZF9c9ves+kYQb9l/bdw4x1bPFYdVp
rAPesQoo9HcSL0vSwQBnApGgoAQhpa5Dz08xpt6ehkgvGN8J17zlU0nMZcPYWWE+
bSu2nQBgHJJWZPx6ttH7pIheQpQkZ/Rgde2g/wai2VsrxJfFwiUSa0LOLgdsy1qZ
DGofJ0x6x5vFS+REg49TAMV3F8x/zUkauqMqtQRvTQUJIjr0FqNn/TkC+HQSz9aF
zUijqRb0RbuOHSq8606ZQQTt21n7PbGysSf+NB0K4CWogqeT8rZluOmRy770eREL
wVVudkK3OkmxG2FeGvGCzZHxpf+AoIZj5fgyducS9Lu6paspUrtd0trm9YjaO5iH
X06tEsuY8cRx3kIczgUcDi89xdP5RrR0W9p0kdz9aCBxYJ+Yg89ExBusiWwT1/5z
OsS67pV7MbaPCG3JfYTdLAjp8ExYjrNgiR9zcHoOced7J9rh6aNreCbSrQtaXAy8
XoRepZQlQiX+MorzunJo4E9qy1kR2NNaGVbHQ5REkPh9ua+sLiN0hDaq1a5LYvDz
N+/QXF15+dOuPJLrKZlwoVWB7hpdZ+yICOovz420DBnRbM24LV3yR7kQa2pqOeoD
KoAuwt9d6aYppWjboVfxdhQLxc7Q1Qth66k+Kyq24C/C3zKoNMEzljUg6GEb7m7q
1VYCTKcGNRclWvf8zJfdadz/Oc399k5nWuMRQS6sHn0l3G2Hpc4j1Rn+I6w4+ukr
n+7sRmN17cQAesjkYJdcY4dmgL05DJcgzc1mqzeZB90OB0opvI2Z5/dgiTurUnRH
mTeKxtYYRjD03YNUDY80+ehbJqHb3+6vaBag0Ljzot+Thydt6klyPN8yNBVvV/iy
tM+lOEBVztimpoh6SU4wLElNsXTWB1yhEd57a8z6Oruw9UFGqCZweXyE7cVJwWfi
U11RyzvNjusztgS93yFTUYF77vAkqq50GQVGXpuOwRjCzz0yLQNxXf8suNu/8PsK
gGC17ma+gfQbtL7lhPtiytFDJ42prJ08thYWghgYvo7vMnpU9w/N6kBsNVcPUykZ
qW+17OOTwfwoBPpE+IdhcwU3dQbXjWg57ecobc7Vmnu88gvAUaeW9ihyPWmT1lcp
88VkymF0xqDTKklNK3MMRhse51m1bEo1dhG4eWMluOXicKWfcFLtzbVxGdjp1O3n
oO+DcefEuck0eznWGia8YJ0Rk+BLPPxS2F5XgCixQXNBVRoO+yQ4osFYxC2rr7cu
DilGqoj25HJy0/QFfXVFucBWlmpDO7bcqqfazqCu2j5yzbWZrpxZKavkpXNAEAUx
NSMHD0aM+bVWXOCpi75e0fS5lymbnESX18/nKpFn+RtERKnohmkdkBeZxHGHlzlj
r50XUSLgWG899eZ4UNcBV2G5gdxlrbBBvv9PUh3gSt+RfkFA50L3rVc+jD4DnzRu
GlT/bCExnhTmo3rok8BUZLvSDN4YI/vz7Q6GfC+H6OFFsrZ/hw1B5T2vshk5qMmw
cSNnXzUFhzd5J7NX9ph4WBrH9cDo/toyS2J2bgfnPV04YqiC/oFEYAIYibT0rCIp
qDLt0M0V1+M7hUKhgkajd1EI/gFZ7HlnW9v+h73gqJ0EjBXaMoXnp/TdJVA94g6M
TMdwo3ryqwAw/mhMARwvqaKT0GSjISH4yHSQz9Ja45KN+zB+yFNFEf6E2IbfyOaY
nRlLI+loM1VGM/Ajqhc0b74ZYkH3hPgfK5Q0mPI5Ts96sMKuW+l5b9v4JUP02s4T
ZKVn9S5NrlEa5hTKWjySG7CBVzjPtnhdddJalawWHurEBkbRquiU5toHQBXeSUO8
JxInpByXi6YZTRfNy4wmrJswUI8okFOiQDbugn6V7D4tihpHl3IJTi1q6Rco2pdv
Z9hfeNZrPwenbbM2+wUR5mlL4x3N7N31iYF29pWzvW5lAl/u7r2A3qM5QqLa6l4S
NudUpMs8ZlYnU1W/ivaV+B/5e5i1pwzp6EjkKwA598zGAmqj6OIGlrslI2iVtXCy
XoLaxrXR4KxJh3TKqcC4mBYeppNrrcI3OWmO9EEvnNPwv12Tj+U1kBlRlJpcLMir
ckD/W+tTEzayASLmOS+DhTiQ5gSQjoJogaIzkSbuVIf9N3o1WkQ8y/UD3hSR7n2Q
gteVZsoLdoYIH9gaAnxWRodDG9FZz90vcoBUcphW40kmDPYuDCg1JI8+QjoS8h0K
s3GjkyeQtyiyIPHn0Ux8OaR1fVM5WIjA4QU8V+6MG7SbbcqaiagbDR+eDz84LvLS
W3bDiiTG7nRe69lGIc2wsVq9XCndxYpN9qwaNHWCwG63p8nrWK97soi7VQrSlhnH
Iw90z8xE6xAJs6eH0YseXbFSB6ZnjOlOHfWGis82flcbyLfo0VGar3qX1MrGuhj7
DmJ3rfNWdP1yv8ab90MvG0cEESWvj+k8znEg486ycXJnoX9IuByckZ+39GJzpNZB
KRrPXhq/cCtORSb1nr1SvVuJtTC8zbT910hZV3WfpiZnt4y8/sWvio/lZo4x0ELf
mf8tn2sMb6ulT/1EZ5opQq/+Im2bCY1oodzqaX80VmfuE9xw+G9HfV0/DkdFm+ED
SQBXR9f74TNJFJy0wk5RvGmA2CMgEOp7rprshdIKX9DMXL6UUJ6Rmq46Udto1nKo
tf4k9EcsJCC6DDZrOWTtBQsK3FF4kkNjY9H2fvY9MCqy84Sb6UUQu49Azx3Yzggx
g5DETmu4Eiem7Gc+FPGOzMeqIf/LIby2v5+FrrRKuo6i1120hny3zyUmHRVihhAh
FZgaRZuJM8U2oejnYYaD22fQU+2Q8YImqbpIa8gsRfMD69JuAUzm+lwWUYwZKXR0
gXY+EEolyhYGCMM2N5f+E1RLJrI+yUvGcaFMXLLfwK4hxnt5vwGXJVX1lv7shTwD
Rhoq1chdLe6iTUqYMJRm36FnY3vYnrU/3nlgq9YYnJ8xlWr6Mo+ZhZANdy+ql5hi
Q5fV7SCvLE68zN2z9uDqdP17bp+bmRejKCXYqOdpzHUNNfmrIuF0gOy+v04mqNk9
MeZiGmW+TcCgQ0e8uhId8RoczrOOyEVrv1qExbk2BhAbDYU4BjLQcg1m16qvS6wM
reM/9QdXr9q3J7j8jPlh0m/KJXA/ALt6XMBuhKB4AkBJfISlmFijpwQGR+kmVv70
TVTxD/oiBiGcK30JLwTeqlULUsTWow+Rl3uWXmfwcK3K8nLv+yhHJfe1sfTNOdw/
mvpVK5AAzYcXrRDjO1kKFDlhWe9A/KiIkBjt8l6o9tAJ8jPQCokXOUb/FHoBHYsj
LwBDAcR6ubxm6AoZVE4qX2p/AxAIpTP0VDxVNE4rtCJ6YqYKAAiinn4tS6UM17WC
IBOAO+9dkKi4q3BFXuxr/O4XeQ7obQ2lTugfXQZdTPLitEz88IpEEBW26YvIgdDx
KHU+6P87PzCKojO76S0pogCjcFKk3q3wt0qicFQszHZ7Nv+yMqIjb61KtZr6KIMh
dfw3iDLBoT1k26ddmFw0eYxQYNwDG24SebWu9WCAdRlIVrPV3+JIkht/NTskJsv1
P7T+K+VLnNjGtr+FYM0+32ALYb+0ZEuWeHLj5aTmcpzbWRDvZThKjoGBa3jXMa5A
Y5aJx0KblucsUIkwGARga4rYIALHeAYrlG3sYjjJddxveyy082sq5Ws3wMNTEniN
pvu9cvP6rDOaJNpcETMNcwO74EWVcau5NgXkx+SOFATLuj8DwVnG+eiQ/Ia5sZ8h
O4j8mxZbHoRnXsjYEP+0UtZ3mFroe4cGjIs/OEHqNa07Rywd6JWcJhXiEKd/SPkO
Pi3KCWMJYl/K/JTPVGriUDmOhkn3+Ta0zkuq4Xs471YmEEwR8x91SLs9Kzqo6IZo
cLZOyQLZhLdSo9yKVnTjqBs28jS2U6lKwJWAdgz2ckG0FqdvAoYdAoJJq6V12TRs
dIxKBXyyS7P60iJ9yXH/Y7lssxWEWDAnasFflHJLt5ToUL7NGshoJktCLyAClNla
VDRBOFYwewiXSJJwe6MdNHJ/fIY9z1t85qWgMHQ27pt/+9DBdO6OP8MCYpwMvzlU
/rpttJvbNDnhd05E8JIqnHJNjmKKyf5edwnBGBJXujo285MqCkRQ3xND4CJLybSH
WkNJgysolCUghlKuXPB3jIa9W9LEnZJJr6nNUuubiFjy/wuVd54A5bOSTxDqt76w
LNGZ4ZiiReo+Y/+0q8nOQ4fmN+sVRQysFCga0nxrBv+NTBlg2SFnd+Yun9/nZJkB
kGg/XiEZtc3W+MIu+oubgwf8wfwpAkJs/iB6HugIlUnV+yuQsIKqHmHuW0JI/4Xm
lOVaXWWaU/7nVrlaEhMd8SFLcLh8YnKyvUWoszGaT2utLrxHlnh6Ly3YW/6xovGH
nyKRt4e5MWpBYHyytV3Yr0FwLNtBs2x7MLdZDHefc0eQFnmL/p82EtlyyvweAb1t
J1Mbfu5f4+7poch7zusbZyqZ6xnwCr+xP9p+BCqlUXaDqOVuUXneDCGwha99snWV
O+sUPq+BJitYvrwUV70fc2CfULfgVXpuDhQB2oM8wsyzsA0OaEQnOGDRsXDUozDK
Xe/2IYiQML1EB2uqVIjTP5jKoBF68Fzvb4Zf4vnPCRA2b4I4JxHlqLy2vqF91hp5
rdW9FiTg7qlYum/gHpuCJwGYEmiJIR9LnxLUYuyMD8ipaJoMqzhkWegs+E9WDSF2
atLEkLw7A597ix4pi+N1PELanl90PIhkKIXiLYsRhyRsL/w5f5AIrb2OfigGMAGC
kzqw17Sz5iw38KSo3jy83GBX7t3sKeFyillcK000op9Tu9M9gwomBxF0WZk2aJg9
hvXZSwbwM9/ai1oGTH03SU/Yk6q71cxOKmyovkvv6KDf/Zgk1rzA8/ZRt8i+Kf4A
csirfF3/tYSiIE98sneCujl/kHNj89/uOcG/LJ2r0YMWu4XE98xMjlKdo93bLOg3
l5zMiXohxoTFYcOUO1haHZhkFOHfo5vMkQdeMhfdme+qPhX4nmQ99vkCK+Zf2HNU
EEnquUs9u0NQGgoA7hyTxyQmtwjFMUk16TQ4M+YsvCRFvS5o10rKZuDyvYUhwlXh
mMNpmFAqUzLGIbJcjB2Lxdm9BAkXtlHojKTRd8BcjujSSeFGdXGs38w0vfwd8uEo
Vw7/tvBeSoR83wdduJx/xwtnjv6xwddN6tJeBvGrPJ+tzlvFnEpeU2xXZX2sdQOj
ZdI9GsFP01sMnQYa5uRSH/bhh+iw3c88opTw7HQY50H/v0b/ixHSJNOQ/4MyxcFw
AedmOgVbP7zOJiAktmBGoXpJncDvLfYoEnKXtgq8wYE36PnddHdNunJMbqd9S755
zDJEb45VyYm9bHrLX5kdhdFIHqO9f97Rov+r8LPn2zVlRazzrPwms77HTo0l/+sQ
HGNyRVPlO1bbKcHXDSLVN0mV/HZUYKEypN+1QpFmr7bOl2mFALkkZvN3phwm7d6y
Wa0ZEFoKYA3hEOLH005mwYE19tizHf6fG/7WTtttmmjyngbnH/qdOAqfYnUuO+qo
naAAhiKqZZ8sypWGdA0qrtffsVdfpPx62SDUIZDymb7cVh0M26kYqCMc12qZhROu
4EghtzVCG3JK9Pbx/aCf4t3iNyY12lhP2Vl4dhWDpgYls4uNEkpB/VJg6K8AHhcv
CyrZJV9R0esBvVIjNh+EX1M0/Af0ewp82qjVY6r7T2BKkGSSbnAWR3smbmQhw60Y
u7onp2auHWb09nM9mz+wfiLiAN/B7l6JagPTTd7r3WWXWb1OKwSwOJE/OKr13Xj+
8FOPGbFoBZEOQlfLJx/uZtKMvOmSGNBKwlRaYScbFPMrMvj/kExyDlkrZtp7DWaz
0SxJPBCWZmPLlpvgsQU4czlcwLMt2m+xG+RetXwPwihidvZT/Km9Ht626snCrxf6
28Qv8gzg2gesW4VOzK9iwhDGaYUlSYOd0PRxlCRMQDBffAuu5d4LFSrbflp2zkC0
775b7Ps0AFCQLNKO9iypcarIS9X5jcGeApswP3YAJ6lAiKXDSAsGPDu6HLzCPLdF
+5lA8TDQI9faRS6VpAo7uD6D9rU4Q7OolESebt/pYV4t72E+QZOy9eLj5vouqJQD
L1/4BsXcX1z3kCUQYp04yM5euynCOQeVr94G4IW3vMFKUn5MEnY6QndIej/6CYEv
AI35b5MLfQjz2qzqphLbrEiFMsAn80Kbn2XFBYZ7rACyVdw5w8Ienf2s5Eqm55q+
ipHdEGoyvjERu4MBnm84T5eL5PdBVMweJuLXIFqkpHRnfEHg/AKp9TaMVn+KALwm
5lAeQ09KA5TCH++9lm1VCk9we1I/nOrPoLjN1KDnRVT/WXspoLnksLaIGPdk8fCw
a9Qe3ox5qay0yxO0Ugnpb/DbCnBl+EWwZ+3ZwGqMqDQXD6RI8H340wUWzJyXFH4d
3JsMwMwVoQNkfOWRwROF9H+M2zYvr0yzIBw4e7KwCnKk7bdWftm+f9xPBa9f4ar5
eCeGM7ecC7QHpJRtF/MlCWOQCdDfJZLbS/B550NDTpRiY9iHYiHWcEyrcJQ6yomt
5aJa4ffE4RqoHcEXkqElJsG0VnB3NLhG8TYZoqGqjCXoXmhe2C8zKHiKJsqwJP92
0f7zB7y4GEElBZywtaJ6dEM7L3Gf/IHneQGvRnE0KNAtKLH/8caYdGVslxcV6vnp
huVMvLH0pAY2nA8b1x9nwqhx/lYs3w5fS1TclA7ajjvFJbFshL8Cscq8X81n3GFv
Cu1jCkbuNMWpkGkVpP5FZMUR/ASTJoa2NYEfNS+6c7BhgBCKquo6p1vlLg4HhLvd
uQDCQpCh1WaoQ80n0CD2zkuVdIxNYqofjitQmlnr/4j9x6IcbYhG/XiCs4td5Q8Y
JTsjQASFtnbhuLP1zCDQm2EnfJQYBme0ivzCKS36PmNVWV9mQ/OiQXoZZdTVyRwV
Axko7hXpK0z5q2welLS+sJeLgDWnLVlMwxlgNCKopf6gimt5TOoLzNGuelr0nkXP
rq7I569EkHtqgmJcDk4m1zS4LKXQNoid3Ek8d1na0EctJcEr51cwog74J7ElrhNQ
Uh93hAHtcSMFgj/i00pAkAUbPdk1pSW78GaGZyGyOt5AOaWwNxMMqb/FhqMcAu8S
cSZaPVA0euNp1Qd+aAXTjeeFfSj+ihBQLNDOkluiYIYkVln7qw4y16lb1EC10T0l
kYY0jwPU/YPIwf/U6zKWZAIObUqAuYttvWkqX9tniSvzaLyJRSZlQydshDft3B4C
NWdHFq/FcEzDs1/ukZZdTaMDxEGeEYUrQHAihJ7CtnO6ImrhF24LF39EYY5pF/cH
QduzuY34RuIYKtex0n4g4SZqpYyNz41CpLpWmrvPQANF8Lfgg4qoiPFfVfUJfrkx
cH6pKKGG8H+1YLNQyeFDNwCgj2c5DxHqGnu4Hrn1vEm9uFpa+FOFKwvH9WJ0Zcx3
BA3dwoTB/ATHXp/dPgrqGEncA9mPbYG75I03KK93fNLKOX0eqDxK2vtcIeBlmRUT
tWqqNALtK3aYG5XCyuTxEeZI2Jacs+1w5WD8Yu28xdg10TXRMSV+x1XGltv3YDum
TDegGDjEMXAXY2aiE3JuJjOduT9i3c94kVFrc9ufU3dGSL4sAGi6i4BInwSfGKTp
kzuaLlynvhKvGdH3N+16L9Jz1DCjPIJv4fkHEMcME4l7VReUv3Fl3wsHQKYSEntW
gFqbiSUrACHDVwL+DkVoDQjmXaBnF3wcXCVxPBoJPX50N2c422JNXM1cFoftxPyJ
34zB4Cq1XF5+SR+8GXsnVZTvyZe2SpQ//KYNCQjmLvquekGn6Eet1YeSWUTQ3zlJ
7xEg34zDm9lr4VmDAduMDEuwRiJYa6N1aX0h94m2Boeuw5soyEpk6Lg7LV1LYIn4
iEnVuYD8uTCxboqZ66NsYFnenNvZOSmKXDgpPmaJfbyJ48vGlRBQrUImKfdKWk5i
0vbQcPDh6zL2mQTfC2V6en/LqTtosoHp8HScubrYC8yZKg8iVDIm6LSaBNurMvsJ
PlxcdcYrOJn/TrQj0LzfD5c6zx5cAqejASsiaQxALQ7A8E1tkOLWyjfy5g0IFT+x
1hRpGGrQeMU1gs3p1Cphp99R3xTrMwFfxTNkhsgfHQu24H2qyd7U/fgck8mttYqc
hTko6xrLnGqB/3UioH9QcbiaxHDTnUNU6xz/8UIlC4psK7+H6RQSGnlygMBBn4Jx
Yk0qaA5sCyslhIYHEkzb50HtCbpufDoKxORVG4n/AfUciRi5InF7NP1eBSUfzM0o
8W41vUm6rAo2LhDH1RZJiE4oFgSU/UWVyve3MqiwosZgc/z7zclOd+3a1wx64jv6
P6H5NU0pwW949v1yOBIfQEnT0Pqm3ILq6GCWFTLvOCJU3XTXf8A0+P13hjPJ03Lr
jYqwlDtfuDybRe13KqaTw2CTdb6X6aAp1oMjPU4zaMnwxuvQIHuy9KEX4Jgokh2e
XBexInnAaAujLeADjZnAFCt/2arharCUrzHx4AkallWNGl4SdLhvCEBSKC8uDZGa
2zFNlwtw778vN1Rq7dX7OdAL5P4f4F1BYEwTW0zsa7kMMnDqJnPHvFEPAy4h2CMf
uLcPRA4K4LZFmby2c6EhHIbKYAQphRS7wJQkRTbz7O5OC7WIFQNnpE163Ep+BLhE
/kO1XBMcAwB38nwTss2IBCwM65azVhJXCGQ7szVOV41Q6gu98GEhbt6D91Ea2Kpe
ksL9ila0jPE6NndOP/gTPQRmvti3qJASn9a0Pz7NSsYCptSSgoo7qFpjVq0eq3tU
MPYQvGZblSi4PSah9V+/7G9Qiix2EPBzN64VzYQCXgmdzbofb/wUyfnAp1+LJRSJ
9mNaF0JsFothP8URbETcugIH/l27o3+0P93YwyBd52LoqAxXd+LsCRqMTve30RvK
PFv8pAmbZqJOzlN/C9+C4NzB8zeikknJaxmg9VN/jRLD8LLteVGzAlt9SORuFErs
F6qLXTUxdFzdbgDawwIeRwHyzxQCw9Hwfsf0v/tQ09GgiuM/q4yQlrJtP+wQ1vAf
KdAxO0mYKTM9TFu+EeEDhrAG0N6hO17BXjl3VK1N26yG66g7pV4q3BydKjBMcPym
mFa+DwYl5GBCUBlGoRjsn2QY/wqIDt+G2xiC4mjdeWZFDTyYv2LKbHiVh6wNRA7N
l47y7cmsIDtj3V0QUy5KDwY+tKcHAv1ileLQC/d+BC3BhDrhIsk2bvHSO3PX3xwj
0N/v7voWKWG6pG8SSbKpoyZrjK5MVpL+KCqQxbXHMve3nh6bAPcR/ucVE8g+mmug
IQ5X2w5vJG1tKvxFuwFYPkLBmqXfurtj5ClwDsfQ6Is9qOrJaBiLraKXRJ6wRQea
FZjXZLjYMS6a1t7YFqOXkirm88JFPQpwXKmAOF2eiZ3+/mt2uxRcyLWUDDk6Ihjy
0X2YE7va4PoYkMDI6pIU0SxuHO24UtSbcyxEzavYEMgmqSw2yWcd5OIFXtbN/4cl
vvJKx4O/aBNNc40S5xZfF55n9a2o2lE5/ebzUfLEjo9AZnXd6Qu4ZPjEHcIJF+Gg
GyaULkMvOx6o0w+Znedk/dEoxlDLa4ReUdICt8NEbXDU5GqefSAZiAywOdWJykzV
GNe+iC600rfRJXqryJtE5JX6795fhXusS7y77EXjxNyYBScmQf/eDOJIo1+HTYML
7XwoS9RRjL/rbERmtkm3B0d6mcv5fjLRwkEXpONF/WU9OAToxNvu2neWTN8Gw5sw
dykrOhCfxf037AU0eFuS8eRAmJ0CVDyLMkzwplwYT6WLYsBaKrPwMvLe1KXD2Ba+
QrUPpTSXGzWTkWby0KVVf2+dJnbiLs0IghAfaqO0BTEZUqFdzvm42H0TBT2W9/dq
dHUt/6JGdl4OCWSbHUUNOkSf9JMhveEHOhU7PFKrI6H6/LZpQ6mpodz6P/c9N7Gx
CCJklJOmr5qPNNyoSICUEFXy6GU8mDAdzKQWnPdWjeLn9Ze3xID/N3O/KTOlnKVE
dGnx4pCufNytobKezJmqMI3E/tfmUJwtW7t5E5gd0FTl1n+dOXiG9TutRHLxRZqB
JVBWgdyZtSoOD309Kddhrt1Ru7MRFc5mFTXfVc7Ps7ihszKJ6SDGlc1j/JQ0Rmd+
PR5w91gS6gzGFVkBVtskNgLjVVcethCyFM9kO7PaPnUk1kdnb/y9a4I16xa9zpxm
bsCu3HLTDcP6WY5Qiaus7ksO3HGi2vGuqbTYdZdHt/Cyg0y0d1ETUW5uY7DUq5qR
EMn/IHtN96rfKtbrkWXcHP5e0b1TgwYzyvsw+3fEx41iNznx8vFF8IBdQBfHsoT1
2i1dT/7nSGy7aAjxvK+jaMJ6CB8hgG0V8NwwWs9Qkw9I49gW4xjh8CpD8Gru+Qmj
D1TzUmvTEpUhK69laRp1/RMdrizxzbIBF5xSTdA22x4FZHxzmKGKM3JykWQ4BUp4
yzVK30DyhI8GV4CsvxOHxk0r54CvId4UBb3CKKXfxDxBkIUwPLUJqLurTo5TKVSv
zDziqWc88Q/U8vtEGPbilYYfPEn5MeUtMV/HQEnLS3NDAEHvsIL0/gMXLf1NwE+x
MoA8DnLbEbMQ+vVe+Ac/BPwU2s3qnG8gHnhxVA85kQMucxACEBwYx3nOP2lOmxDq
Odj2VGSRMED9Zndz7xwLf5yHIUjikVXDU1/c67aMQowIGNpDCw7IHqfj9OmWJIja
CljijuF2R6dXoFZDlJZMFLBJ1G7tqxLDVCLWjwCY1+c83xsa2h4YqsJWidcByqcZ
Y54J1qvV3X6ZVboHQ7BcLpQrM1gt0h4UtNAJMRhD/M/ABfpnDiW0TJOelKDI28mh
MM52aPtUzSlmlKXiYrGF/mck9L6OBh/XIUPj4O+1wMg/blM/OA7DUG5wuFlV/NMz
MFWevM5Alt/sfMGHEQ/APDftmfRApGJRcoOVECSJVe15P9I3/T51HQGzKrPstqvs
z1+LxgDXinmXtKXYSPiqzv4QmIBMatJIoyDSEe1Ibu/KgBTib8wGCvHBvfUxaAz4
lAmlwgGmL+7V0BpeN4Qd+ku9yEXknd8j8/1+UWSh2ioubQ10vCjeitlNyQG62qgU
Ekkrz8dAzXlljgIa+BQG3zQuMNxmdym9CYJZm4JOt7Ez8adAuxOVdil5/Bi1PiwN
fnynzNoH2TTXBqD2jvW5jGg+II669gnghtoeWzdjfYGdR2mJf4pk5LJ3kvL8ETgz
y5LivAkZ6arrfiUzsVluAvuf5G2JmsTvD3yUBJ5CLIDmrKF0QMkErS0RrVB5jhFd
jSIfKjKVfspowcw208M1bZpd0gu22/P2bEkRV43enROhBOExJgOnL031nUYdfypX
kLQCWo4Qvi+n2OEmri9NNbu13y33ICTREAvbzB8Z8lhUxhIM+OOtOrqVe9yMxjF/
gLPKxn1fZC3T2ZtvFi0VCPAXQO64WNuIrvjhNAqCSvb2mm9V/RUNgGnoG0ZgzLeo
HQaKGy+x0n4TRQk6DaYH6gw99cLwxpyYgxAHIMJGWSNo1r5jRRZjGnCrnoKQCqmz
DSfQI9lTnis+cnJehYmYxCoXUPX+cNJZwFr4G6mZZrDN2+vtNFBaa6l9CC9vIsYg
uL5RTQtENek2U555m+1CFYNdMsXL+O4ABPJZY4Ng/0s8VKXqKio/FMU3NJhgWAOX
hb9TxMm2UHUPWYMgihQNbNsU9psfeeW7sISJYUTQ8shBv79J0GJRJ+5UMZ3bxLJ1
NGkyqs0R6g6Axz7Y4qpw0MTzp7PUyOSRzyJWJFejwMqSj/Rg+2LmL4LUQjxgs30Q
hTwpkOHGEeEukZKwNipyLtoqFQgB3vvQcW9nMemKyIcfceRQG3B/Bn5+L7uymoLi
KHpH0RqM61OZFlZuAB3bwh0Bt4KIws6Afkb7DbcT/14ji/ZIcJ0G8FSJp1CXlNKn
wEfcPkCZ2KY9unBBjtrU2Q+dCfAgB72Nslpo3is+WuXkS+dcNP+KBHDWhmZ2wwNt
XfGmJ2nlTSik/t7vDM/chrnSK3A9ZO+H9sdvw5Z+l2tD2+7eMrTIjk1kchzXYK2K
5o4Dji0tSrNxaGaj02npl8u6PVZO/gnRyI5sC+92LuUg4v1oREYMG1N77Hjupvh6
PIJCv85BSvHDC+9GqeqeNbq3pSJUvbfP2AR4C7RwEqSHiicKVBR92lyLmRY+1zRt
SkDkokOihG+7UWPkARDzfb35WGB8MzX3JUinNmvaKdhCnXQ3eD/0Acu+MvSC9Fuj
rWFif2Hfs/j+YMT6/jeitkZxo4vluWXePjxnPPLu4ZukDHTMhF7eh5om0y1wsB/e
JE+r/Ev2l4vAYq5RHCJEsSlZ83AGKoaTR/N92Dm+Mq5qMeT1uvH3zReG0jd/DMf1
RRjN3Wzp5pQX8GbwSMwmroEByo+azh2MB/ZaMxC5ANHqihecsau/UyR3VD6kuSi5
50VUYk564WtH2gQ1Ms9Re0DrgjRvIXq0YpbDeJ5jyyHxh/a4gHfdICwmGV4QnxNK
F3ExXXSQumbDovSIZmCcogg295HKFLGQrRHKEbpRvRxHR1AQSftuAtxhVcad19xH
d0DcMLBAbWnLRxeBvJls2XuvIpxmM9wbh1N+nlibVAuZvYwI1LIK1Ka9ejQiJI19
UA1DTfoP79RcNvNvQYhDpZEkuguJUDCEGxLNcDwaqy8/hIAvQp3x0NJu9SYIYpC3
xWBxvdJkI3SBj94HvpCW6pG8OyqIG7EVlZT6MZKv/wED1j8x9GXh+pgBiDyDxt8m
7UTy5MyTlqiCLRC+Xlw13pgGrgomH2tvhlZ8ZRby3pXDaJd4v2T5E7txehvs+C3X
FG4a3NzecEP1y5wTfa2ckDB+Qpjz3tz7HLd4bFaQ9FDdmn0jKhX2FQ7kNjTeF75m
wOtZ1WSfTq+4wvacArGNpIHRYKDq3y/r7ga955qho3U2IOhg6ZNqBYeWVbAY2I+X
nLAT3ARjlVmsNiH+RAZp1eXGa1ptjEMG9sdFgeflB0GIRWaa+TwUX0slJByyuypq
Jp3rLQQ4o1krFchsIznWzW/pc79KFrnLeub0e1KjFfaFIiuzC09RZwOYIH2cKa45
6XMLg7km7fbgQNgsTHdzT60Zy/vvefY+zjl+WgFBHVHgaoGrYKSeDZKr2l2p92ax
B8lRAteog/eplilVHzPY23D5Jx/pO8UTMbWy61CVOPDTGJ6mhSmWdxRkIpi+MNUo
AIXzL9MPqOOftvnTwmnIHLpUe2YLfjX80xBJ/+WyhhN/Lq7o9OtuAo2kjCgFgqrN
FKZ5FN/kKKsporQWQnV1assWG/XY2/mNFKrRQAL1CX6XQ6dleCEp1sEQoD7KgnR9
oFhLJ117tsD8VNA9VPQvPtGMout1zNl3MvEt23FJ3txc7/BnMctVAciskDyVBGI6
aBwR9ucSoipiLENzGCx1oaC/jwfoCLPobnZ6JkC6b4ISjmZVIOiG/U+wLfYkDlgF
UpaviMH4mrni9dXCbTVL5ZYKZcg/tuSffzIFclD2P8xUacuOW8ohYzHOmEjob08h
jxUr1nL7hgu/a8g6scSObc5IEW9WBfNX8afJ94lZOxeYFevkpY8CRB95wUiHFzAk
9SrY4lt3QYqExXaZhQTWtQJHgsDu+KP/xE+zZ3tYjW0xpypNFWz3v+XQmWaiHA7d
4rYQvRdP9VRQxzgNAbqTM2HQRqeZDdv23aGJavh1vS25SPuuouYBB4RyHv2ShYs8
SolALTeXesu6anvxWM9sAnQ1+Mfihss37tAzkGvRIRI4tMHdRJbzbW6FV5gU1lrA
VxTAMZmywXjXUm9CeP5mSm8VlJBNuR6mJ1On/ckC7NG73hvbog6Dcc8wMEp1nVAd
1XmwnlnB+ptufOkK+zfzJr7QZNvOmaXnjyYwJkhXTG59XjKCEKs5FfKbhrG9P7T3
POAedDxTCzYgMWZJrM2cMeqV0W+aNoN/ENFrBqkQQHNXIb3saBqL2ZUI0SH5Oq3Q
MFE1I+5KlfslbziIq8y84OUNFOTSIqSVhi93YpTTkE9OmARMZWi0s+0ivkCHWypf
U4Tpnal++efhDjupOAslMh4JRpB14hJ2qhD4YvkUht8igFjDRpYQ7tjehHErXXEQ
+0mPoN2HIC/vVZOJO5TXXffTC4GAytQHVNhKEasKTRYzNhPnlYWBwe3uNyfGRIsH
uN77AM2fZi+lt7/OSeFJHDNf+rXl+LmvfiuJrbZrQchWoL/T2a3W8+zbWbQ9khVz
QORSkmzXutDvzJ6yFcC3WoQO3lBQvchxTPUkPSr/cyctpcjJvsIVZs3iPSebohqm
ka7cG3Up9InTm8jmZEnMBu0TJWv5C3WurdyMJ7YcaWzP0I9m1IgGAaUclABaqfeD
CgMBPtYnDkUbOYzdod7cRNf3mQ/jtMbzPYCYOnQKpzPxcfsdH1iHygD0QXUZr0wc
QFIuimpEb6frRzmAy8kOkEXd3bvW8sptyuwpZfuYdnt1QQFeKWvj26o+bFo7fINN
mMdqEV4mU9flXbhNqoGpPokCqmvUAjx5jfSH3cfRNXlsb0TIc2RENpDBbmFxJQB3
awbMImkquR9DoM3zfBr1thyY0Qn40E7Epnb+w7SCmzU8col+Dj72gB+hlOhjOz5E
TFhDLVGD3II4jXrGmuLUEcSXto76BtSAKAOnmB8YVd3Xau6a3yXbHU/LHdqy4TAA
NjquEkqeqSMStevHb3hpyH+rRd/0LUjuqD3zCfENno89k0PQXnAu8lJzrGkTGEly
DgaBWptiXS2xl/wkWvuKxdOIPZ/iUGtGol/eN/CmqKrfxRSpj7a/kdG86IKHBLQV
RVS6xFMhkf1+ajLCl1RkQokPXaqvZmibyT6pMdeaYZCCAhhu+VQf1uexABbJrPXv
DJ528UOvuIIbKwUXPzRbk6B8CjrirszViUTvt2pJ9YsCRKc73WNrCC9NMdArex1W
mLjPhwP85dWoZBxh80JEY2mDsfi6ZzUKHhas9oilwbynECKyjdxmBEYxc/HBsATx
Uj+wK6JJeLLuJCN6AY4OAwBNzoCj9rJ9lQDo+rNtgcz++MHrjPT2CMBE0RKujq42
dtZvAF15at0jkS5fpBbVHorTEpKY52RcR3PBwyOEUOpHpZUbkOfItRsCzYtpq+/a
X06vbSQm/BGqoBy9NUk+gh7Eh5XGSgg5Z2ItafKfRjw5Paatddr17fczj8rdJ31b
BhawR3+OSHxhOMG/ICoEJi+hc1BmQP7ropFWAbdf9+4ey1NLVpce8XM6Z0FU1bCj
d1qBt8ufQe9NYZMKBGVGO8cR3xVpPuLnhZLgjJRVk11Wjhh2LHC3z7y3Y4hh+VyX
n4sg9AcP3stWdaKHpKS7A6rXwC/zkIGJl6Z/hz0Umij/Bcp1VXwrh29aKz3b16y5
TU65RkJ8TXFnaO99DrrELdoBJ+3eRDc5ccz6h+c/roWpo8OYg1p1akRdt7AuMivB
CMFfdNNTTnSYxcEcspYUndQU2Dk+gBDI8jUtsngxUdtTVaO4v+i1pbOfBP3GScUi
p4NSN3NsGn+/qm2n9rRpNuEegY8vk3TRxcd2/BH/yzI9lvadOUnP/cvSceJZQcgL
9ECroxsBfWZT3MlX6zz8HcJkb7Qt2EZjU1yOiXJXQ2d/mUZjVnWXYGME22cPynb9
rAz9T912FhbAobuuFf4Y5BAzUXWnnm5186hS4PI3aVBrrrlRp1nuhCGlYRyXxzX3
mhoWGjsFsw+bnLzYQ8xab1F82EA+qD4mmuM1P9nkXedEjfC4lpHjkrvMz3Fvao/p
NlX5mhwlKy2AJ0XhSse4k7uMMlYBNOFZ/prjCxcFtBgH+ecPzrjns+MBtTRMCB9B
VzmLhWKjIvkIfslfCmLGJa3qY/1yPRYkBKi9fqcFZv/LKwgu2jhBgw4VK8+jc4up
RiF+K4q8laUP2Y/9WoOpEAe0gCahBJvtVRDbQbbsb7hFhSqPfKLYkaNN+KbfR58b
1GsOGDnOmpLrCG7RbNHT0wueYJO39Z3zkpWZpaJGb38LDbdYDKUzwYiK7cjZxUwR
Bhnkt8TB5CaVmzdeTgwt/V/hHTlehLrEzA/mD1EuLtJ1nrrZLggWWJ/1Lwa19TEo
7q4LF3lBUQc6aBkdkKmFWGh/WrJE/lZb8SYnxa+nlrMr6JEbTErjpYgi3abparFY
mymppeXe3H43qT3H5QTI6TeekoaNzlP44ppDSmPt/8thNzLgYEj8nr7bsMAmv99J
KsoBFTIDCfWC4sbq9rUtvoRCPmTqOhiOFJxJ+U4CokTGtGpZV1LyemMtaTe9AWvN
zckx5QVMW/zCdMkfLgy7IbvAZXWlznvwsg9mM0S2NisHwWeof/gdld/z0ImXlCt2
FstY6++iAdcf217tt6lTh8aC8QGIlz1YjuoPGxWzSAyVaHmkhIEhlSn+z9dHbD7Q
zofwsR+dDaJ80gPAbcNMaIDJGezVfdoRAl7XV570Z5M3pygzhtmo5JTqRbNwaQAe
agFGmviZnqpZ6741V7O5spd+LoX3R/okAzDci9tacBMVNnNzBQazu33ElfRorxsS
UCsF2vpDPQu/H5lPJaHAHVzaE4vOAFrxzWIWg4SFxHU1KyFSyiS5YdbtIKEc0XAx
9wBiBedGC5n+FtjYUmnTtrM4BdZOGiyBcncAFjtZ7PZUc03+4CAKbwtyV2CPbKAM
nd9OLqee0Vgh6lTuf7S4a5pK3nFNBS5x4pYpdhlie9PsDh5eon4wTeew7ncgul7/
QCrpf2glU6i8USQgrtqC9tMYG7UDV6/Adea2kXs7APVMo4jTqhiOY865L5OgwgHP
BXG/878GCdRovNDhm/EH666SogXNxIflBByyWLCXLoUkKSHsEAhJDTpAKkCXJ6Mj
tJexmiEOaBQos+g51MRutyvC5m3hFaypwtTVz+w9eK3hSCOvEdf3NuUUDXOFSFGE
HN3B8giMiYZNju8JSW/fmeSWaxX7S3lBEUOWzw6rwOBlNyvh62U2Ho1vwWxpoClR
KquaX1s74DHltu/DVQ72oQ28NQhs5Uhe74cyTny0VSI6wOxiLB9RrH5xbKETFKrg
ehe8sYO1GWvTwICjiuKYIzKSNqdG91w3+iCmr+v4Y20NAz+STI3AdaPA9TIZdd1H
pyFZ/X2fYZCHAfZjcf/zcq2KbVCExgV9WyHmYBtnNNECDeX/Ia5MQGgRYEfiheLn
m2ZQlinmQkr0YN83EJ4hBcB/y196sUlSZlG2aGKW/C0m4zV3Ux5ZVxVSTslyVOCH
mssViXWZ4rYLuB3T87bYqilrotoFUBmjWbQUGdyhBiJ1Z6sCv/5cJOIhO2Hem5NO
WUGxVRTSxfs9BxcpQd3FoSwAHsU+bcyczjNfT9kSKPxE4nlBTKQgL8+WaqdhNh0P
Vlj7WvlmckE3gTb/eILc4IsQebSgyFg7Z1nkPP017f6u0+MeAmJ2eVagCDJ8FXlH
O5WoXL7bQay28jT2sLhhStgJwCYqOpOEft+7XRKhy8v4/cjqP8wkBIWVimwqX7AO
6DEq3YVTJs0YKa/9ZuUtLzy3mfTLpVKseXXc0X3ozlrrwHtwLezNb3MZGt+ZqgPm
PNNKI/v4jJzQWO4srmSTA7FQOEMenHFybf2EZT2xP02QY6ReMlUNapuiFev32GaG
nvO8ybhhpfbUn1bmAfrJs1HlzHdmnGfZdVqD6qjHn6vUsP50niSucWUiXkpWjDUW
/xs8kOQnkvlxtBGhtqLzgG4n6l+Cbg5PEf/phM8wA+eSpjr6AcOcBOWEnAPsnswk
iDG4oxFmVxVcsa3JhCOX/25VmApDJCR1tEopw0D80EgLq20sVHdNyq66CXZQXmNf
sS+VZ+vhJ2Zh2BzFE23iTy2UQZIzd1dgVhiLQBZ3lawZBj1dVnL686NPFKSF0IZ7
Bik9f5lUcTj4dWaI4+Mhz53GuMFlNMtnhRmB88OZbZAtZe0ahheOE2BBsWUXrH2z
H4Kv5VmurhNSDxiqJUY8XVb+3gRyXE2GGLnjg5DIQPCYsP5VMlA+ToS3iL5XaBbE
AeyN6Bjm4rdd/uSPfzS9wVW7sRRNUfGAh0P25PAjz6Mt+jmV4ROK7xcsZyT5nUmd
i+//1QX/mq/GggeZc8Y2+d8NjzxEe8pa3e2y5JNB5ZA6/4TQdlsBWp4qjzFW7np0
wH0ut2xwfwlUZo0ZOUmen97MlXGhrLZdDjodmbIY2vXTrd+gOc8jdVCwBW1Nn2J2
4v+fM8CxQvP8W8rxYDMVDUgyA6o3azqZvMmTncvMSbWA7aPgiVpqC3fx67uMz5Z+
Z4FJ2LCtrWb6oikInsCvU1SQ+rD6325m7YKlQ3V7I9e/Ss+kq6kMO9U15hbduU7r
jN4Pz/2b/7yStxYjeriNyaaWTVsjP3M9c3Xd8DraNTVC3FqXdnr1BP5tSpLvgVzm
fvVHwpAmAid19SG+ec8L6wJ4EGYdA2XaHEGyGQOW0Zi3TFteOo7Rd71rssDQ3pha
I55BJE2LLCG/BBfyr3lUiS67e1KGvFXhP0twCY2hMwinlJ2550Tx+ND4ueQgbtew
720kFWJdU1Mag93YZ49V6mGcNebbeNF+Xvryu78LhL36ZR/ta0b16cO2ivTUavMu
WxBEtmTZbPEjpOZl68JBWBOtYuh+iSUY4rMURE0Z/XU+/wKT8IC1AP4vHg1bKmFV
oTijESuzP1smEC/IW0r05EMF9onCVU1NNmbBaLlDv9WtM1R14BSBz1tJs7eyszEY
TysbKyfN5zuim6Zk8QLqtzYfHP2BjD0+6tNZoLi7s4AH5TiBOdnfdpWf8SYib2LB
rnG2npplrZI1TIKxSgV1CiRFUNupow7zwTvyaPAV+0rdwfalIlJiL30ctbwtn5M7
mQoy06jnk4ryJmineOdtwjNCENWecnnlYtpgXnhx1YDurvImBp++2LBUeZWCrLoS
33Hx53vpZdUoi5zfCdJZe6/qYBok0sxa/vfidJcFybvXLrmlibPHupaBE/xPPIKL
soA/Dm9dPihJsmaFZgCBeKY5Rz6XYNIiziqCDNuGxzXklFkXO0VVoLfd/3BpmTsk
R/dUfViKUReTpZ+976OB3toSsTU2iu4MKI5JpLJwm8Q0P8o0PjmyEEU9H4KKbufp
ZJxEW3DivpM21Dz354OkQdD91uEUtr8lTN748WSRQEGMzJF4oLTRrlXeNx6X1FWn
bebZ7iRZsfU0vxFNd7emODLRlS118YGgPynKRa3x0zumpfhYqI0xyqKMc850RU5Y
xWGWVf6K1f2Q7/3EfnucCvgCVeI1M3jP2/bwds3++vyYEUl459L0K8kqLYeRWltI
dx9sVyCc2S5I+xCfS1pcsLtj8ivud45CdoJGM1i3tX3ufFMPeJb23xcbMCxVU/LD
2YZ0spBqLxr4ADX7RB7sK06Cdbq2U74+CRoRX9YYOnZNxvylE6TS28Yc5gJ10v8A
3prj5mqRoI8JtuTGyQ8M8ErK5f6hs3SLVA382ujYDa4Y+OZFJLv8GgNshtBsKJaU
o4H/T8xW3zM5rr1VRCjyHM4KkfkQUiHzsXZyqpvw/B2fI80PERH9AtgrLwSIk1LQ
13tgM/wPiyyYpS034SZAU9KXE9vQdbONpnofsYFjapyLO245gEuzumLHStU0iovE
Ce/fqg/9+LxdLPyyFYTw1HVhy1zPXXOsfvHIUjna5S9xQ7R5nTWJpsi6pcVo6ocq
D5/qxuZQj1p3xNVMlLCkb8HBcqQa4nvh52LpMeHmgxPiqXSUI+MCfToaBhCl/Y+l
CWUpCeBRcwfbMSt0JLNzUj6Zz/BcKWZqcS8Aestrg3ddTMlFTdpGzHMxuaggnJ/E
pxUJVE6MwNRolFFToM9MyvzfVSX+P2WnEnXB8WyV8marhhtMwYNJlGlgNN9mejHb
cctF1r1tzCJQEqqZu732fXDcShh8QohAyUNtB7FlKz1dlVRdx2ePqUwwbxWHNVzT
BlQYL4/MqPAs2iVChEY/k3XOjLOWE1G6Gyi79Qkfy/iESeYKsuinjwUkY7N4ZXjs
fdJED3xu+WJu+erstXaKSRbLy1MzdW5Edc4YquYt9rSqoNbXhwnTIY9NlQQ9Glqp
xIU9J/8zeJyAviHcQ1cjHY+0OluOz14YyTBwyB2RxNy7Z6Byf8ju88/vp8mI5ggf
lrXCTnfAhBYMKCN+Wx+/cxM+w8p6PFa9c65CkdJsrTgl1BeA6vzbnRBRsy14cQYR
BdsdVCQ6Nqwmf5PtbTVPWnIojgFuNSibQK6rlMWOLxCc0u/9MMIXs3WN2+K+WPyN
Fj+tHGt8QAx7EEKhGuI2enQaSoaKJkih2lxqNNNxjEkdukjuiu3guFwAeqY63Lj0
93LcgbPgmJc3RsBGs6xbMBKY+0LDm2UfPSx3qNAduW7PTcZvmmjlt6srsbzSid/R
l3OVph4fM4+X/FihQWyVeXPWv7ohD9fVrpEQ8k0FVKvvrLISXQbHYR33QtIjZnHu
X8yA71OXZgoZB5SNkXVpcr2ZrysLHek8uXVDkGDc5iiiKuPw8PgYBF0K4ulkyedR
s9CfIRAPGiNGWT36SFzrqheKS4oaTn3q3/kdJaZay2mbo0uWYSMJkB0S8YFSq9f7
e7Q6WDLHWX2yE/XaWrbIJJIds+YrAdrY47l9VMGIKmMXrHnVNT/wA08PdGvvy6tk
5KSmQmhyHJbQ9srTVw+aifmGqOQvV7Ar0SXZ/rhnBybE7v6NFsC/bxbbyl+5bIA7
R5v5/3zogKzDmmNNAR1J0uZlHZYjTWtenAjjcbNY/A8ITFGBHChtDrytAAiaC82c
LXAinEyhn4HhSxGPCv4l17xnoxfCeTttga+cGiSO1/5LvSxHgfaMzAX61cYOs3of
4l7eU8b0j+Psofny/EykSUV5iKGxOQtIrUd3C9z+3fbc7iacJNrLPrc/TrMvvlzl
mYEcnQWPRlIrEywcmXeVcb297OvLcObrHYQje6wNa2jV4yI9DHoEQqzHQStL4kNp
wxFncKO0fuVO1ltAwHBBXrXX5VRNT/gLVYuyyVtymaSMytkJ1FG2Fkpkln25EYS3
irlSS18RcwKW4yGqB8EPvp2zWqus0jPGWwivyoULT3VabMQf3dnllE1FAU/JRWOu
OUFGR07Vh7ri0/qy8skW8htUOuPdt8JXHP4TCp/EbVBp3xQO1N4pcaxVhb+MiFUF
YdXocQsuir3OjOOba2mCTXTTX9bdPuwKQQp76fUCm7b0Tvlqcj9t5Liy0XBw4Ilf
wi08HxThnO+73GMm7dQfTR6s4BZLVqMUKOilbKtA3eyahvR8HHdZO28HL7UUCYmW
/5EqgGGyh+ll4e9WLH+Ks0wY5VaqAvtGclgGFOoHH6ZjKAjnrxexCCwz4hNDH5+M
/PLYu4ZjfGTfgPtDtzOuXMt8vZxMp/7jTtQbRJdUrxRLrX+h6C0aACPaEVSKpYOT
yJ8FSq/vKFaMG+O9hDFWSH7o+luc9GbJhI8brhAIWaSwXnm8dWlZnpWJYHe7La9v
WQEYNB9dXZnUQvqXHkK/CKlS7oXADEXWyagBhgZCCAsmDFRUccaX7JjXm3p00dgW
bQMxEa5pF+qcgtous8MS/0gla0FXQeCPKg9XBD9ktI5kkanQyDVX4/mL7lnQVJ1x
l2+e+rw46NxX/aHGgSAA/DRR+9AQdNYqx58bhZ+PojmZdo6BTAfU5OoqzBfq+U7+
pFTpbP7KTXS8G64SjcFEYeLAqmnpdps94vGu45KfZh6aKWqt/3r+bwDnRvSagscj
aWuWe01iUUF87tyllxy7G+e2B6eoPrq90opEuHPqpcAZG0Dug8/KR62tzSsZnEe8
yVJpUcRrBbj/vfpSrKrp4wopkjSUD3wc0Yz1zZ91h64nzkJkLmijXhWBSR5eSDFd
0eBmsNTMLYwC+sGCVd32oMZN28eYNLbx9ZQFLnkBs1ubYgefYpjFz+EsYn85Y2m0
jNa9BTyiWH/KNpSzqH9dtnwy4eprOPHtxz6u3p2khqR3x9DYaWoxepHY1goICe+O
MhR56EWjZorPWJ8MXajwjbqh9gdgZjFCCdVeflF3dnJIOpy6jU+RP+V/Tye7+aXV
/H9SFb8H+DYGPz4tBe8yJI/1Ev0x/djfy7O9dcmbIh1fAa7npd9BxEoXxDg+bXfJ
V7kylYZ8ob6QLzHPXijLsZvkLq3U9DWkc1FqFpngno8wucw4HZ+wMpFPqnKxZkd9
Fjua/kJbGl8JerozdythZPkTdjqg13eMGzGjFygRFvDVpW9yscqVanLvck6Z3/X+
M8qYXPRdP3UvekeSZStPQTgWvSY4GS1PQpylw424s+G4PadzGu7/rSWTO/fjTczj
B4JJRTIh1nwRXGhhIJpUwtaT9ImTpLOhoU3OSBgMICjHZwkn8sjbIxfimSqouDOC
OZEEQlV61CGNccfP+6lVGCO63FR2rYVeHkSabr/A2PV37ANMxhDGb0WNYOvKWfnM
X01XwvcgU+zcAIQkAhtAuh6GTGAZdJ1JKopBSfT3TVRniwXTu6F7BBdz5Er4m9eG
aSGhwtbbkgnnxXP1zjFUeoO3EDWS8x8bCgIf19W0+znzjYCCUWjw47bHsksYHLKR
VZ+EQ8GXgSt7ftvAKLN2byU1wQ7BE24HivsM1vqf2SGcRI0CpuujOiR7LrdDArIp
SV+7ddJm6fzoFI3NjOuaUXmRnUt9Hp3qJRVV+LidUQT2Olt6RUYILGHDd1HHpPwO
wZfrjBQZ/5XYL6kAKKlqrkQUobDpK7TGWA0w35aH4rmALCKGYdMFXFDOyT8PsvUL
17qvjrUIRT2VheK4e1XYJ9RI01s2gYs9rLtUhu0ut0W2veypNwjxGIrT6vKG6RLM
1ZTXe2BuMiEP2aqYyK6tKaa+wi3fZmRBWAVkyZ1eDUEV4kGmcTsaKn5UX9MJqH4i
uqYXW5RuVcNyYx773dS1zDKSmQz+KRx//+LGAPZlIIBfH73L6WUXHxesk3G6DlHP
5o+4gHiCmJW2/UDATPi1MVQiQsir3DKMXIJeRrG9u6qLdzZikI7X0nXNM37qUabU
nc5g5Uc1D+tanDpRTnTrxmbSvZ6tpKDbPBY0IZ3cskJK5EMCKsN61Y/1/3AYf8ID
8iW1ZalgBGxAxN+VfMFfBWPGk474X3mW6HsUMiL/jjZogvOG7lc7qisoUVVlqeRO
NySBUr+q6nnIk6LICvryz8OIV/Ai/9Kug5zRXCofoa5+tTkqsTBVIO7uYm36MOYE
gWWnHnvM0t1SPKPJNedhKwps6EYGNITdva3QutCrl3P16tXxWlu4NoSs6Km64hB+
zieJQgG6aVNbIyIhPF7dXJEyTNgAOARt8RAOwuUYxPhbDalixmrW25zfotExRr6t
SEzlsiWh+WjNJrYtlr9nIrrZsMQHYZlWdQ4uUEGvfHTTMUrA14LWSKHkouitc/aK
SC4nO0XL2nOhA8kvXymQt+MGU3P+0D1w1KSklKh5kQTVMPokEH/TQEz6K0lCl1zs
au/LKC0wBpsn6ub8N8AcQq9SYnMt4xcp87gEBV95I2XnvylUbLSzkdppTpBSEVvr
Jn7mGAyeO1waDFes9z3FX4sVrUBksdmOg/Mo0WOZhh9QGNd9UXb96j16AOf1rHKi
uHQgG6k/cFfF8TLqv69iYEdiMKkFGjZhtjR94fCM3Q7hyzeiSRw5zhtLDlby5i8r
3CDZnpeZfRkiPYNm8yHjTMOw+2csIUDKSxKy09bdyh3VtIdODRNJUrLV31zpxnNg
ykUshnGvvTnie5sGPn8JI013f6f+h3/rN5T/ZNrqrmSSnhxafWyN+7cFm7Ib7oCB
yxmkfmXmoL/5i70phDY5XJLoMdduar046M73Xr4aY2CMdcGWx6VKhUdDm/uXM+dq
syGn8FTsbV2D+SjbWV1Co47kgvroprNSRmXSBvKAJcn0F+lDXk79jvL4hb2ZkhyC
V4T41Gf0cfbntWHRFTd8rJ6rBiUQO0R0S5fH3nwytAY/UtO2MEBdjpzg7m73915W
HK+VRQDS6epiiqzebR68qDc1EDSWqsqgtZAdVCfpTREpwc4ePXJVGYd5p1DJcdQQ
ykUnfaU1G052K3o3hqTWwHGEV1XfVV5oX6sbEz+PAiE/k8QqqAmzQi/l43JREQTM
WFUh54tLZnWzLlE0zrbqYtrdF0y6xxQP8kHj283RaJINCg4F1BvdhTdimIfKQaCs
b0HMD9pEkNdDqIRGZ9i+Ezfn9Xkc5+4JsdgbvUn/TgzJ4KADSVHIxxj/lfbR0Vjd
LJgF28XmOF7934I89dsoozxeOQNoLL5CxSgpWVzkWqv67eAclpLMC3Z2eshl5Dd+
MbqTu1sHSfDD6m2mHtCm9YEIti/oCqCzv54D13/6PTv8VDJRWywqAjB712UWT7Kr
Msm8fZ10nfcVKufgX2Ds4fEhqAhiXDEd3+coddFRtmHVkU4RNIXYnViRuE8jfLWq
RrG+4b/M4+tqcMspwPWUkff46ge7zWq+mO2uMYsSZLpv0s8+WAJXWSa3polK1AbZ
T4UabLNcBoFHDXwThBm00lODv4k/P21Mr0fRcVEUyWhFzN0bNCSFwSEtucvzpAp0
V6pywW3zDconV9fuZ6WvLi9DWt00qpvcd9UUNMbqkNSfj/UtGsz7lwNaSu4+q5yX
K2SYq6pHXc30aBXkmYczT/Hn0zcdMr7y/ld17lXE8/mrml3919riAb2ZLsJqGdJn
B9ekcWPxauPVmOOtKfjDp8srRQhROBFRxa32y+OzBKFvi3j8OxVAONrGL/cqz2WT
PkulPq/L42JP0c58mfZjnU+Ab/zXLm+rDx3Yif/FCcGebym0cmSrUo6CXXtW9E1C
s5d+1RZ2eTonoLf230giEPnQe/XZDdH/aDPOBl/EaMN1HuQmBjKg0PxdTWj6YOPP
AoWpt8juZUrVnFVDQ5xatmT3M/mR8QUJz2Br9ehdlYv64cUMWd3A7VYzjvGcymf5
iCzj9ctg4WL3fzuk1gNRK5iqEmm2ZD2nei2sI2KuMeS/HmaZ+poquNjtdF23aSGW
qVw2akTlWR2yJ9MVB/bCdFo+Y838W15qt/HANhGwIteXM/zIyYwBKiALio6Nc8Du
PcTIdEV0+oo2aKAridYE1ZRCnUyLEU80e+fD6Wh1CRlxLc2uetp0rJBVFvbeldL4
xl7JGpHFMDQAJyZ6I0zU14JhP2rrgBYL1lxvwPItoD/v7u8MR6qb5YALf4ttMAxD
F9fdhe7/hR3NlwHaF+BhY2xN5NdQu4MpbCuolYoBaum/b+CqMpoIFvLIAIjaa+ZA
HVEqsI2HFtaP6IxSBTP8Hggjx8s9MyHQNSYPPtc1y9J/xitAqsd4DYt3D3u+rM03
+RtjkXeUCkrhCtRecULh1xglb4Gt8wEnuy0/hHU7XrbXb+G1sid54LmpN9EkC1YR
Sn+S64NYub9WeIWl7wMll3oPHOOn9gakIGE3YBxuPU3Eezrf73VYAMY/OaBYMQsF
AwEcVFkhp3NHFv8culzfd4aXFXS0kvj8NdiUcketzUHFPbtQCpq9qB4WmAajD1Vg
g4CWfnD6HLbvw8YuYw/sAvkmo7pBconaa8fNkMT/RuGDHmVaMtoEJxLEnQXrMCK/
lQAakvezU3B2Mi2vvlhmGEhTEYsEPGkyMXA0Uz/yUW0qQmwsY1xtjm+m/g5xZxWL
Pprr0HjmO36JREXGoLXtg5kMNVywzkplPA178EAmeJ/A53gMwrdgqel3xlT0bHwE
Yvz/gwzBdQgnYdUtK0LfY0+TwztNwywv5MDCuXRuV9ugUh/4ch6DEs8KBH43jfIX
qgLgRrJ85b7d04d7ZLTM+cWi9V6LBMt7OzMBlde+nQvBUyqdDdEtzuymGsR+t/Cw
Pvr2jQIl8jqlSdoK5fJGT9bBDeuq234ZDnnWqp/vs9t2P+/2DsL03xAVsPGu1qNu
dqZXdoKVjjVyyBuvjwc/nHnh5XsycTpPDAj20PQvjOpNkcVW2qKP0/OBlLzChSUf
MW2KkSD/QM4MzjzBGZgmi2DrRrSAxVHGkekZlIPWZVwQD/Lw2WPPhcBMla64PZF7
ytJ4OY8KZ2+e+ewM7bvd9Ftqq7/Z5/WY5ScStiER48QIOo91h398iCYlK5lPf2bg
vro/LCPC79fzbTlwiFpYJMKqmCXwz4Z3NyjsToSBdnGIcnvpPVJGVjpkIGHkIKVy
/pztWDkZwSvLOGKA9924GH3NUMOcszqaX0z9CS2JEHTSqKaYZiT72SwHtOSD5lA7
AkpKN5mSH10xUBNfhTp9wOgfGtWI85uVOSMNPmPbR5L/thB3yB5g74lBbXhMRP6e
i9pQ3fzdJk8Zok0+0HjZ2rxrMOhDDD2SF5CQzhFIZQHxWMJZw6xwCH0DdFSIybt4
6gGOROliaWPobEbWFQtwq1DiSq8Tcth+q27PggISO0HK3Cv+JtX8G7TOGhIfsjfr
`pragma protect end_protected
