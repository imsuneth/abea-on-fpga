// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:44 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i9V92eBv468SIXLLHDTMkNxm2qHRgqa4veWExPs6zXs5PXS1FrCHnCiT3Zes2+p8
b3hBgMzNKFItbgF2EDriZ0HHobDy90NlLMunCqrGEp9pLufUWv/9auJ4C5gi7DKw
vSFsNUm8OEODj/1w4QuhoGoEhGStqgBam87z7UazU5s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
g4OjilMbVVm4yBBx+SP2KOv0YPoqFLc4iy9puoWbaeeVIG8EaCO2tjuME6Nhf8HU
pvgtKzS0dLSMKSbZZyXlB3qtYx6bFZO732hIPHGxdWKRfOx1WJQ97M3jK7Q8aOgJ
OvLE8eLgzPJgudu3mVV61Ku8n7TUvo2+Tzn9DBTWtbrUyOg2EEF+4AfWbnKZL05j
TOrz7C661Zbic14LbqjJtUZj1FH0Oem2d7a9bPyfPzvOUsWjR1+en2BOrqu5NeV/
EA/gRnjES629qCV98KdYImfghwO9MW2OfhlY8fiAl8JsaHGturA1/eDgG1QwHQqq
vjHFGQHgFiMwD4JelfJaW/JxuKvZ++1wWbTlsaWO4BrNSbPHj3ryxuQZNvihruSX
yb6N50m/QyqadliEcDOmY9AsQVyRe6Ee/cVSTBj3SKys4YKF0cUCSrWRsXWjFgmB
uqcu14OUHhcby0ndCYKoUxiouzw0KRfrUflbpSi7Aq67Bzy49fLKxipC7mRG1cDU
9yahpr77UVKlDc1+s3AcJMiUO0QjbaKYN8m0lv9/PlG/dYQnzoNqQO/f960ouS0P
fzsquS3+kYdINH4G2gar6io8LKdCzM04M9V9YKtpBojB/qXaaElp72Ys/QEtIBs1
ask9nIi2cY2xMvThTDbGUWKpE/7Xe+Ioio7yf+KV1fY78PDg+6toCfi84uxHuQxL
TP0qmcx7XXihlnLSZpuX2AU8q6Se4BoubGvyqWRbXy6AFLWtWBw6c4Mxlb8vicI0
ONYdW7OATlTtitfCkarkowpNmWBFKMtgyLi7KZArbCmDMRhjj+C3rdMPRj5Dqvdf
/EJ+o7jOeTsnjFuaKMrmRwYRVC2a0ax0KzOIgMpftWtEIUEn56oSlva9/fmIZdkY
0V8xqLk4iwK645MC+Fs3URr+mU+KG7NvtlCEzr/SUbcGwiNlclopMQp0oLVI5kkZ
wHhPnWkKJREh85knSO1e6kE6K/t09JwJdluHacVT2Pc5sdjTQV+IKh7IyBl+TP1D
Y6UxKwh9cNWvt8gzbOHcHh23mThmodAidIqBmL8bfSaFPw0MFI1bCxplwbcrrrKA
Yt6NICg+BJza2b3Icrb/zy0Vfs+QNIROMgUf0t84YHLw/fK/hXkF0qBgTMfuAuBx
ju0nXj2EryctRqgN+p4NWRDP9KJYFX6U+LeM10lfm/q7GOtokdktM9I+P647kggx
chwmo57vIxmM6xqqJOmzY7ez1BISrexbQlkZlXPTeNmqWNUdCxCQWlRI/u+yfMkT
hI+BZS7uidKjn/xZYGgsVyT9kAOVnYH0pKlAeFsamLN7kiy6fCWeg5DF5TzPmO9M
l94s1R6XfAW31GU6EHOsUbTI4/0KuOzd0sOOm/coclh8V/Y/vpC1gHiKNoUvZN8z
Wn+HkFloiswPdLwFyfGFmjaVjqURDnkMKZM7pr3yy/w159QnvpnRMjo0Jnr37SFw
d0Frg2YusCgvrQlZ4imnbfV5PHvOKES60tDOTqy2dsHkC9VsLGybKrc4X5YssRnj
hqU76hFQ4xBfy+JaJOSH2ynQGyX+NqZ+ASolhpUsPbuujSa2ItgPoqnOLY1tW8cB
l1zuo3LK+0fHxPKf1vdVfV6DXiBfC4FnCFIzGU4HATYnYdM2+tolatFjHYQKNUIe
Yt1tTFRD/+aM1Kq/+MhJ8RgCC7Sn4Z/jyUbMJ34pmfyW0Sc8noIlXVNGUMYabdvO
1uCigr+UBQpesfeqlFlU/Ej/IJoYS7Rta+jbFjt0lc13tq+N9YpT5nWTfRDY0LXi
s/wlTSb/2UKa3Tt3FdflqgvnFpShzYk6GL7caSwP0cy1BDwprREx0Av8WcVJ1Kp5
HLWZhEoMBmyH89ZDJk7gZYlXNi0M4C8jFxizDJqyu5VZd68ato9uNjd5IHK97LEt
3C9e4MraFdaqlOnr1S+oE6CG0PWTpHOAoT+HNOGE/M0fauZd6p7IbxqlDfgQjrce
INN55ZKh189XsiCGJiINuckNVhXlqBpEB6A81UKMHx/GRyScMuoeGm5BE3dwVvsj
BLBgQ5zZIyZJWKhs8vEE2tsgegJKjQSMB5QW+Bzk5lMLnec9NOEeOvRCUxPa70hN
MFkHx6jVL75hwhRn2RJQIA1aTZ3u1ZQYnpGLn4NbifT4YGimIbXRTBZctz9FrmPs
qpBVWsRNWYnLDMuUuQEee8BSj0d/f+aDCgXRemCXEba57T0MRdYUvvPUN4kBFKSS
Pm9V+mxrmn4wR6HjC+c4uroZBbh6yB5lFupkR5tV86il64bqLlywWgQ4HsxdUBa8
CWiR7ri4JboO10krqqblzDfh0N2gf91rFRnjB31Y9ng5oS2OHiqd1lc6nEu84CVA
JgxNCmrnWdVb1pqx9scf6snDWNWWCTqRSnvAYnyI7VW3FYZ7BxWUIigp9rRQ9VgE
sa91fG+ZyR6PaAcuHa+cRhPnYTGFzTkEvhiXrQ2cLjTfbbPKIU2bnH35A7PkzGb+
t3gokZxakVTJd7oPL0W4LV00pyNpey1AGC+Sm5RkWUmwYWEePK+535N3sm3y4rC3
17/gqox+HBbG1TzHaOz2IkNEzjYnEOM9Mx3uzEnmtx55tCH1viydUtGHmLRxr6P3
jLHs8Kv9n/MKO6EHWz78aZE8/v9o05HOdoe0k0STVNaJm6+UBfwlPa+H0Qgkiloi
Xryz4ylIluWZI+Egkm5VGY25Ryl1FthL3AgIBvuKGPcnstx3AZio5cCpSGZRMie9
AFlPvJv0WJRCnxRoVZwfRKnQ+bmNNBhzxmHw2tChnT3T7LHbeJggMNV+Dm5qJZwQ
LMkTu6pFP2+RDit+2OOMGROiDKJ7/VB2fhRFyqlDXh5dvPs7NCvAFEMsY9J3pkhK
kcyMQW9FXXeHumsCuaSlUeCr+43YLIuvLiFTKS15Mp9emsigilw5+7NpAMtuOaBl
/iAhb/G5pt2THueYPER4paeI9ITtWv+8Og1ChW5Xdb6HLSefUNp6cQZ6Uuo4id+t
8Yqt85ydnCRjG8oSgbqBPKrYemvJmvrsUG11KHzqL8sxw1ndynauGUiAZvc/7wzj
Qu/zqKinw7DXpil69woNpglhwkMdqioFU6WhaP89kjPar5/d36c8F/W9yYbedVsx
2Zfn/xpiaAWnfC36qF2nPC/Z9RAXxLFNMXQI9dvD4L+ioyPj6rSqA0ucNmZEc46o
TxZGtTyBf3rvZsXgzr1tk1ukfc7Y19ijm8SLuOfPI9oETN2RUrTX+3rvzg7WO1Pg
xKgQncN1+P7xwvRrnpKMmPU3GspxPqPYiPDBBHFDR6twaRZmo3RfloNk9mJoTYhF
30+pd2LLlu9COvB0qjY4E1kbjfpj7nSsQNJUVU6R2G7jTVtxc4kSlTHCd2M98aN2
q1uMx2BfyzKwv7BCCgVjJHefNKFkssZDDUpx1hW7ZPGKG//KpfEbH/W81ReDgfr/
NwEyhDvkqMVm8cVBqSF3LoNhfstv3q7SSEr7c1/MF3qdVEWA67zll6RaI1OTZ7zt
LfKwB+T4W+4y8SGEZULVnEJIbbTA1bW81ik8vqCNG1gj+iaik3y694kiSd7AiTC+
V+KjnyAGRXL8G5chhZBNueiQPdCNkQ9ZV9ElRyNzzCxrXNgaK6s4ZJVeBH3UYr+u
fCQdkC2JxMSw13FySse+s6Dq/idL+nJsBY0SPVcEs7Jpnv9MT010eYcVjQvHRFV+
ZwCC2DA8FuCS3MIOBNH1ELPc+sqcSEacyJrhAQ0yKJrfxuGO1jYw7+dkmeND1zND
4PbMP3miYyhqpoaFITXJYoUz1/dc/ixLcmhxUMvZY9h2ngO+7jruE/Q2eaaG9dg6
OWMLVTfgL3SbVEKxiOEJ+6eFUunCelozO4409Jrvfz6UKId1tAOVrX1e36i4SQFs
wnDmdBrim7TYdDTA9wz+Ais9d4MtYkEsKUMZqMuuz8gfIR21+4im2j0wLIpuN1Tu
WE1kaWv/GRWPVJKNkD4X0n5FTPCLS9Z8fBdBMBx+8+zNxkD4jh8iSrNudcG61i/i
tP3EBtkvMYkmVyDuwxDsGemYrWY5bXgJXCHIzqK2HvGkEzuOXxmncu7n64ifxiFh
04HBrHuEYDQ2MBeCPW4uEq2itPnQrWFK7HVtgg1bSPmPrY7+t0WIERMyeoJo8fqo
IP/vO4Rjp2DshWC854f70P2K0+Wbs2jttCJY/DGzRQpyD6bUUYNGO34yghjA4fnJ
tEVpufuNhoIkrVHJe8VU7P3rBwzLzE5xoaGCpA+bHaOxDma00gL6oTKmgVq7PCFs
omfc03sFnM9v6m3Oxv7t68R8QmSY0zXoudJoFH+Gsn/1ZEE3ifxhfok9I13OIuIa
OvQmq1VWAxW9DuJPRxJrYoiEyv4YC3w4obNP1kbX2O+IVaJ3stBCSnaLQlQAanKV
R0gxmzh9Zqeo0FacSOBecsQpl5iG0xXPrIJKPyqcMcwY9D7u9L5LwsyXAtA1hdcm
Ysx1GkWEWGNvhpl3b5b60ijCXKbqcCVYPM1Yb8uJVja1CnsugUD3m9WnoH1xnGrb
asMPt3OzFCeim8+bY2bKLjNpBklyLSXit9yfZU6O9T2QExI2bRnVDBOiEEeEIOiX
TokmgaH9wZ1y4OAlnBrY5z7vqSVqU9o0fsPaUPOLxB1BsZZnL5oaPEV/qkQnRMrR
MGLuFapIVjuj4CXaWM/DCq8o1S3JQxCPbi9vGedZD2/6L7fSRtshNRHKPGVbthrd
2shEI6mJ2Vg86ZD6c09GPrw2AuNR5fm1BBwUMhK9zfQ9RS90VuxHhx+9ZK2WzV0/
K6VvikAOUJcEbt37mdY6Uuv1AxQIv8n2eQRN3eDBLJkfp8AFXZWRkmDLZD+geY10
an8w48k3/YgASYUhmRP6futeHBEux/bhIbFw7q6ebzCsToAjdsA0g3Wuz0AdUk6M
wvOwPHdFIzo3JgA4L5UfHOjVli/MwecKNw12W6fd83v+l0ttTgxsgPrl7PfsZ872
sQ0DqSmsVIJqscBpd6UUlRGLfnos4eT7x6mSpEQURos1CQS7og9QARislZl5AbRe
q9WpwrEMbSlOUtbQcrhDQrfy6biC6AB+jKtHwOYFehyPUaDrZZqGmJZrEx8GM+KU
19c9C7QPg8bjlpEogJV/MM35lHYvD2rzrdrbAXWTx5g8QY1B6E1yD2GTD/lhWf/l
TAi2KngKtzblt9sRsjFbmembMKOpf0/CRGNuJKO2dzH52LZRnsPdhhznxGnSa9ur
SZvRQCeb4UTrWE3J1kSE0hQu381BSuR2o0WQ+o1Uz5YpMil3IXCLDKuildzBSjcq
/q745MUE7ea0hXu1Enp5KeFppRJuKhgOdda0PZk/hmD5OODt7hgbnNlOIehNHYhX
cqArmR3r6eVOUSudDWcn3xm6fLCIvmL0SQUMOlEZAv4qRFiZliz96XbhPxGLqM53
ufkexjnPuAxdLM+kbnJJLW4yVEjyMnAuyeq3DCHG+0GKbhWzD1+cXA/x5Qtwpax+
YoFUBScHwoSLTElTZkz/vSGumnYZUe9iKe4F8QDkAPiIOIQn65GvqxdR2dLs85Is
jaU+7ql4vyZ/1Ot89JFEkNV2RgrvH68/PeOBOyDUWiRelrBSD4rhSUvs0ba8cJnl
o7hamTzHhHMZhr6w/dJeVs2AC0YEYVag03xQLV3zCkWvZ0CVjS7c3CLuMxBkVdBc
1fesoy2zO8J0bl6s/coTjzxEa1SmKgrEfw5G/92MLL4ybtqpE/3xoxIJeH3M5AMN
qHkX4w83SIK/gaCxOlYu2E+psMgg1T3S1zFasJbV0g0YFz8Re4ENOq9YVnckGgsR
LCyaxL01BCLf/wcLqfqAVCWRCp0LnoKCE4LLLodWSGoV1i2jtNvoQ4iKNCUDvvov
oFljk1nChYhmQD8LgcPTH3csNrNUyeOT6BlLvwLErtw6+8y9M9jFDWl4qEXIcoqQ
Trr5wJueYipSjLYNPAmQa+FKj4dirJl+Og8D61ZszhhO0DqgWOnj1c5xA2q2X4PO
/2PGHfY/kGwocsEIBV3JSL2LxVPVCRzGx7b2B2sJN3D5/d/5Skxw21ABPj9fIfKP
dxflbQL0Ac7vJEGaZkmX+onXKbP9nZzzqVY3oowSo1BEcop8wrvr+1Vqd2jqbmIZ
1QVo4Jo5zpqxxAOVN9LB/0m/dPL2MxS64kzXJyfmzKJUhz6jisWc3cqUTBFkdz4j
IYoHNzfFaNzZ8l8i69CB5leZOPeox1ttx4cNyKznbWb9cfJbOtoSrhCcY5s+a1dL
ZLfbP57PmsqX9h029FH0zS2tqQ920AmrIdKYw/GhwLDzr2u2okG5xyKv+jXkedB7
iZDfkqjwIdmZnKpYF7pz+SPxEoak7WTroeRbPd+O7YRzuZ1sh1babRvdOjQ8SmuG
kNswO5oFnDEeBEE9EVdaNvqgbL8hvY98mebWLoJDuah5NJP5iMKQiuXOgDjaLZZT
EiewB5uGMFhMkq5xjhlXybCxQt1+wANWFSNuTGUIGm9ObXzr2+ULJm+wTtVNSd9W
u7xzF1j+M6egzY7xBj3FuoJAqPWiZGnvHaCVQC72d5KlE4MPU2zQlSpRdlq4l9tL
H8aH7oN+GJ4L5oN4IYqARDgHH8R2jjVGtPim8oV3S7BdLdfMtyUF6WhGPO7O7kVg
OxXdcXB1IJvsTM02ZqHEvT9rwSRk45u+fvvzHffApy1cskOrgm1jegPB9Ti8/OSN
6OKAMo6ZtUKpyz2UMUHjOyr3zhA9kF5Nm7ChKl7BokaXhcJawCvWucH7ht0zEPtj
5/RZ5lsj1JHadVQf4iKxqStrcvGrimGF5otSi6vZYAjPheZv0bOasSt8Kt8DI/+S
9XVt+Q6BN6S5KIX3ZwJrHcciU8s6l+jzSG04N7h6kPrE9gx12lAhAB/C+OrYKQTS
UerSRdeNWrNCmbygduIWYq6IAUZiMzb5fhFJCCz3JbvXNsYtY7HPaHKKLMlKkJsz
OHkZQdIO9G+et5YCMyRE3/UKrlntpz/BT0PK+RmPuAeZwHKoEdvdZh7NtDt/M8vY
eb8Rwq2HZ5KnxRM8F3vLTQoNQZv/tABnOf2BCd4cEec77YWVR2bd4FwbnSAAosRN
vemx9cP5HPIF2Wiki7EEgu78WNsu7duxjuHZ14Ws2//RLA5TM6fc6QRbuE+qZ/Wh
3iXw/jlnpWSJuHe1Jl6VkiRHfhdMOhy6sgg5c2DB+DWg0Yh3fZtdcJxnzlHMRsHl
75/oS9iZDnbN5Qmz/265SlQDLmxfHbfaKuRFHunsSPWQ+NFAtDrmseM47bLEARcG
PrLreH67+Y3Des6YfRWLtnQFlDKutiGbZ3R8Md1ePgUQlB9VejSMHioBLB+USFVp
5gbAsFgk8QAzSANOvYLkbq30+SxDJQgDKPKuSCxAYWALOMN/WkOxq5lEnNImlQuE
05ux/5xHMAqJ925eGzTZybeHszykIlsP4Edx5h6d/zbmMsE3zVlygo1pVQqwAWwg
OWGcA8XOAlQ5IcjeKmyI9EAmXaxN6n32NOfULHSkFl0seLlZ5hp7lc7irMoajJAU
y00zWCUNjSzRevvlkc0bhGSGtUIB8jtOjFmOhkd0JRFEOEK33pKf/e+jM6WcEX+/
`pragma protect end_protected
