// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 03:56:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KTA9xQO7qwYyFIQcLUFxMUsMQL72jjZZoRi+FDqV+AY5im3LaJGuAANkavU3Lvdu
p9ADlexXF115BP5k4v5L2fwhzXaMb1b4uhquMHIN+zHpYHFvLY9DLN+SRK1vgmyG
XJ8Po0lhQZAxGB49BP/0sMsmb1tbc8l8dNArzyGJiNQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
mcnL9+t3hhZaVvwVoqlZtpRYqnvprRTvaHjBXizQbsF96+GGRD+hkR+vWLfHlmqX
u/2tL3tpZX+TtYHaOxtoahM6ZwXxeEj9b4AE9SudsOUHD9cFXyERlpWMUrshYkqx
qJ7LhQG8jTkY1WbxSE5cL21emkMsPSXJjMwPO5t5HUPz+A5kuNRLjWAvEQxKvfaN
4VadNLubuOWszZuvSRmvaguYYdrqZiykJXynCx6+1CbO5ybF0OGKSuKK4LgAHW4/
XB7KiuvLwhTn6vGFCWeaq+RfLDEbDzMUFWAkJzSu54kIHb1uVJc87+wQdK25Q/yV
T/Cs10tpBwFa4yFt7krqcSuTV+Rxh73whWCjpILiWqDuDl3MdTNZJhQU/EK0A3a/
eWtq7O7XIO5cRxxgKgMjd4Ye5/KVZxo+h1TIBOfkELUaJgM04B9j93AOEx0DcvLj
97t/JJhYoCVr5hwQtHrNLcDJSX7Hi0FfMXxGoXFIttyfmmj9+Tcig3fhvMiquO2w
GdhN/kS2AvGjBc/ZwuzDWKuqSOb2xkZYYXCgnZWN7m3z65zaenFczhw9/u3Sp1um
PpWh5p8WX7+FO9KOlJ8yv65ByXpAioR/lBJcAgN3WeeVTjAxJYrrYcQ9mrseVMsO
TWL25KWbsk8zVf1POD/oYa7Fa8LqHtF12C/+u+kLc8X7dLHt3tqr1TGg1eU9q/ea
U5fz3g80JFrPwxWWEL/ukYEAZ3skHaYiOeRpsoLuVCLue2Ygwt68YRHdLcnEQX9k
/AWJK1qpQLpPjcRpCTtKUJ/Wt/qNxj17GUP3TpmVirQVCE2ylCw5vi1rw0xEVOEL
QySEsDN6Lp5tqods5Qj8O0EfO40cnEmhI/2+iGE6ec8Uu2ccnanC+uokW9MfPh1B
HH/hXjAMgj+OMDbOxSe0Rq9wj/3kqSXPosefkV94zWYergdxNbkB6+mH+OQNUZ13
1lcrjhOieTFtiNTV0/q9hVRMA3aGkCGJZ3au8+e4Ujk+MOWexbP7hE3Jy0tgH0vD
qYRCC9HWLC+7XpiYGCuqU6GK37pW++b4JJMePuF+OiIdgF0qfrk4Tg45nXcXJXE7
/5QarA0iwBo1GeKPMeAp7YJTSrhR8uo2qH5IQwteZHRp+QvoV5zj2ayrCcc+U2V1
skQDZh0YSrzOpjR8n7kRBpi2wsbO0iDsf6lw7ztghGUkMR3aOZptlxAj7q23UJv3
CoknsFpPIYdAOy9ef+w0zzI+LpqpHfOYboAJNDwZv0EWkJ3CP6Vr0UXAferTiBLH
dwxEF2q8jjkvHRt/8dlOHiDviA1yogVVsJ3EOJpJBKQ3+2o7sz5zXW2/Nbelwr+Q
DoFDUgu0/lq5jQQvUbCJhienrZOfTHkoImhgBvyFzfobJBHWxBCiMJCAI0hPeysE
qa6F4mZCVExBZ+LVZhp16lZL/Dh7eOclc03ihJ3PtSOc4WwBVcgt4cZ49D10N1WQ
HuoaTd0H9Bj4EBbLUaemmlnWQH/b5rJLN+o2TvI3NIKe+e8G2YYjgP4kEW8+Nt7C
aXqAAzh7kMrWrJkztw2UKnyjWGei8vIVABujQt2l3VduzU93fepDxVKgyPOFRx2G
nJgzIDtu86bMKXPm8idf5AoA5nuB/SK/21zswo8kW3UHJvWxOXBMV6p6CVMxdqYl
mrrnoMJjz9TMOF99TlgdBxUbZL9PR4BDdpIIYleCT58yQ0JoXHyNtAS3Zsbog0FW
E50vcMKR8eh6i9AlV4wzKyL0rLFB+kZLRNGGKNN/vXAGj7bqSk3OnTdIEycSxPhE
2Fl20w+LJS9LainTKsDgB+Bm60n6w19rUIKKeSz6bcRBNR68vC44mIcoJLYekNwB
fyNlH4J9yK6Ahijlr+sRbj1cK1iEHHurhSHNHQJrX2CdPzdsnfqWwvYjicIZmlku
/UGxar9GMVP1s7KqKRbMBQXwIvOzyBPFzvUamcPhbsTK+NS8oelQFPWatFZlgTPW
KboI/lW2PAS4fMqyh42mhsDWXnUzGws5MHtr0QjugqPtBHph5I+e4phbsgJkIfZ8
td8jpQE1qkJWJpFA2AD3DpctVhl2pGBl67YJYNh+3YzW952TqOYZqu7LV7iJgAgq
Ek/ALkKASPLbSvkYADgVQoNPrKPCAkiO0eMjuL2HaquCkcXs0/pldeolHW0kKFY2
Ha7ihY/fHN9Z2+2+gCUDbpQ9FQ0QVCcJzuTWtRUz8v83u12XPvs8m72fJRwrr425
yW8mOFG2zhGkEoyGdqcZDRVn45iuMIEw4/HcYWc5cdhJbHGfbT6X20EzkfpFm3A0
oDOmThYHqZliZW6Z24aTwMsE5IqzQupT9K8GEhpWXBjt2KTpQE05F1osNXaK85h0
r/9I6KkPXu3O8iZZtQhTu4qbOKGNSE6SYay/kNAyRW/dnrgUQFSNDvcBuNIB42sU
ZatIQYaM8Z9ADdNPdzept/GsBeDrtsgWeiztjuLJQbZQ0w1vkfQeDFEkWlj/ahTy
nBwEYXRVrmgx0w7TNqOTVTXYOwUWmu2E46So0Udim2sxCbtXpS5rTcuE1AcI5kD+
izG2fijfggjFxsdftXVc4Tit18pxZK0GW4Xa5BiiIeBc1SoQoo/toSPoKnz3miGR
OPdMU/C3O9Ahiu3RyduTgE/Jdwj//15nyBtC3Gi96BJFiuFE85R8CR6pQCDGvQqQ
jdtnMAGVKKCtcYLoOOUFyLnWT977ZNL6xlIn1hC41ImjDH5NLbuyCcduBVQCly1O
FvInVKL6xV7/izY8ehPNIKeQ4WY9idtYqm3k0gyDaeDm9nqkYMAxHBmhCvvdwdmK
lsH4u5Jw3h9C0OUKLLRamo03IEmj/Zqj6ZljzgFdfeSbnfnjeoBnHG015H/kS9dF
twrZEE4fAfRmn91KfOQMfIh9akLM2ge5D0HiuVugEJzt9+ENTiT6Z0y4rWBWK94d
ecpxGc7BRzh7O2A6ekGq/Be3zeWt8+ka300vp0z6DikzxUcUY/AprbrqnmhfED4v
1fjl0TvmYFHN2TSHIkrX9Vky8sCcDP7HQJnVHDpZ1VIyCaK4nqCih2GL27ZlDbny
SLNPfBc/zqNmpqlKvdNlAJW1gk3bFbBiJMN9tDrITu2xGf1KBq8N1gk5pA4s2ixU
jUTNsuv9E+omMzcaOXxDW80NMYd5dAMmMGHSyk/q6wPU0MbspTSWriSH8OwulsZT
WAHV7FRRODbtmP+m2hvfLi2TroO9CIfFa9RNaiaumiN7zYlBHHNLwbOvY4iI0TM2
oX3i+L6GyLVNGGwvT1R331T0/aRd26rT0YnpgwhYE+uEIh20+Cq+CFZxHmQoEmhq
OCok9VXzgJzY6yvyMmYWJbTr2B0E1AvqoB89Jj3fo6j2uPwGbSPr/j31M3F5omcP
xNryAweMFuduCUhxF0JgWaCZUDonZv/H7fAC9J0cDchLYYsjVqtdiBdVSfZd6eHL
KH1I+6TK+iQuqCtJiDCiMMomwiWb0yP+mfkR+Pu4mnyj0uy2NTWM4v8NBj1atK6W
jgcVAyMZIw6pQx3WuhUhGSFkERhz3GS8dz5Red/vB7ZGb3fR33CSJN8StIyfbLIw
sda2OzA3Qlps/CCg/iLuveDpwIHaUOdKLmjl/EIoW/UuWxkZgAmhQwVgzRgP1Qcp
C0EGT9WvUhqXAPGIvJMvUzyKZKQci1LQZ5yEEAM2XxcyFguCWZ9s30Hf0qAY+laD
gkF+IcySdKGHb0Pprhft7cI9+ZdNV2rQiT8UYN5iBF5yVOOXYJiXf/dlHVi+jhKF
bcQhfgu50A2MOJF05GJWLkWVwTTXxLnfKh8hxojHbiKfJ9oGLOxAuIXyVNoFjNZ6
YNjMbPtGqH6HszOyGTbqfjZek6d8IWNKJcPn3is3IsSNXKvWr+SouW92BInsggdB
F2EGbArSmTVFJAGks7qZEUvhO7G8fk5CQ8kEQqTOFrWtfbhZiQ4WHZBHxPQMf2rY
D2N/yLJVHnO+ihoPT+BifEnld0QBK6bN/Dmxq5SSBGJQxI12a8rwDS+dB/Q0ghS0
iQXhg+USMI+wgXDCVUSK+FgYDVD6/LLITK/+sTUuFQ6XbB6qboS9LnGG4W0RqmQF
QD3b5cFAC5COtsZ1A6K0U5RiISIJFGX3emy7vm4iI7DY7lMYzeLDvNBKP5ZGFZRP
qO+sjjvOVRqUiNHhVFgJIK8qIV17fkwiYWPCGyu4yfCCDnbeip5y7U9iOAWrcJ5l
h5RlNdt+eAP07O7vaS8JRb1VlI3QLn98uki0ociasM2VjFoxmpSg0HFjMGFzXhQ+
lFU81ctB1RMJ6QGZ11voGrrTV+zN+XkDxq757oIpGu5a9ifJ4GutTIE0q3PQlBfj
gNb9tqVxUqqNSBuRsri0KwQEfi1muT7UvcEIwZ4XoatZxk1obH35wZrcvOFyFj7Z
t9KR69xXMcXFdyAuRScRDxBP0NDwfI4+YxeMaRwmWeunodAk82JJy9TYwSm6tV1g
Ld4SJ3xvCa3VzL5uoQPJMPu4040BA/FZjBcOhDOM7V51vbt9E6GmsnbNUGXFr1JW
V4uuhRppiNIGC9wElPzXEz3yhuFQ719ik6g6BOaDKnxn6E7zx1hUtrxJSbJ8S66J
T8pzA87931VD2vzKoGUn/9ogOLIxsHz2ux+VufULXTtYUC+NpR1CRYJadBbYdUdW
BbItsdbaRJ1C8VuoWTxAt5jV8reasSRDPRnNc3xMRO5Bb+ScQMDYDhTF1bLr6Df3
NY9r9H1W0kelO8bJDnivyZPRRZtM1d+3SJRiqALls6pSKe1k8uF/X2PE5+Qae3RH
j5eXhQa/KWdmjXQnqril9EBHTRJ8wUlqSELQNF0MRY105g5DvR9ILuvH/bAOy5FO
eld0TLK7gpkI1coZSz5uJq8/NDX/8JkSldLyrANNqzue3hUdpRMUGT5fLc4zCvSY
XKNIBVXPCPf70cc36LSIGgAPLCiLrXU9Mo3uK/n/7CRBQPRPYpOxwOdQkOwO1eGH
VNrHL49N2PHz0R0wzxzsAks9ZHpEp9wLYBBXbrnRFz9ceFAt3md2wWs6uR+ruOCV
AIhE796bIEeN9NnqvpEbRv0ep5bmru8KV9QXtKtvfHEX3XbpVhLk6l9JA3MhpcEG
rJgypoDGDowM2LXUCvENke6pPFgeVTbjsA6MLm7SVNL71bB8X/clMPc0xX8ECC4W
Cx6EFHkJHIy3WhhNMf2nmo3fnbtT1RvsTXDnlui/G26E0DxsBp6wwJZL9zG7TuFx
fu3dluBgOhvgAx9Q/qpS7rcvLQUEe8vxs+muJb3UUqU0270g/Bw3S9ryN9KiizV6
JMPtsRWMTr+liCtpqrn2yi+HIRoLUYsWz69RK/tzcgYMwZeNJkKK1EVTe4FSwTLd
w+SlN22HQj2a9Zw/p6Z+gF4BkIuT3YpiQ+h2qFVbc4BRK866PbLrlyNLM58QEshn
W8nvY8KlmQq4WU/6KocvefyfT6N3WT3j8SVvQfLQQ1PB5REBLybL2ptxBEybDQ6V
ldYQSi0kKGMlzaIpz+oEaLuRBJKXbuDXfTFa1XiHARhAVOFbTGVhMvs4i1kfA/Y1
Id7sDr8aQOsJgVT3roQY2WsBHaXS5rmwxLOCFkFsU3bASS7WqpKiY5CA9J7S4hgv
jqER4pDG8t9pmJ4ZNn1rYRgzFd9AWyKr38P/1uBTntUbpBPZXZfWcBPJZV0ORRfv
nClH4U1676+RlYOyFb69Q/mRpMBIBJQ+dsTbep/23K1ZjJmEdW2pn3ob7j3zQYmz
z+8j+Q7rl5qgczP335MDx1gB4dRuQX2Wy2DmVKYRCMN/0+/VDl58tTfXjKS10NAn
GFUCkQUUfOCWOc5rOAIUGMBWqIWWUMra7CYWaC2uhtejOdd5kafYBBxWax1bQPRr
f2s0WzZVADvPUKbqDKligjZB0vXFVU+ty91KkPM3ZNGzPFCpw+A7eCum4WA1uvka
B1Wk2OIWAg/8LiPnLOjodHhW/6Hj+tknt+elANDu5NtDdShXUmeYA/lwR9EzFI9c
AwNiJ/XJBin9C61zqBJkpSpGIwp0T3j8BROptcURjRDY72jFseX2A9ZWqJV+BjrN
hoRFROcbPiT+qToxXzd2khshTk6vvPfWh/yQaWgDY4qLDAm/B+WBg4iyCTGoVOYD
KtnzG/vX9gL8+rNsK8T/wkamjTfm1SkY4KxxWxgb88XpJEX2xDTrjcCCWk53EjYf
S29VmufWPpQZQ/VI4oDpsMJaTj5Qo1VoP1BUEA2Jfz+Kf6pFZfiIWl6GW6MXAZ3Y
8yfvdH4ZBnberBrQZwS3IZP3fQF2OB74irXaXauniKZDC73sI5VICKDW+Gimo04S
C5HmuN09mS/M0X+Ncayb+VrsIOr90/roUER006jDzZho2t+fPzrn5eW060QLjX7s
aZFFK4iekY769Xcmh72WejCJcJBCVS4xUm1jHzgdaPLy9xHEOlbmXsYN96imtldI
PZ01lSstqPe8xcU0bd7DjfOaM3Jd2WgxEI7q6v4opHj7nYKUcvNkdHiw+h+59sAb
BBgCmUjPECzaonF186P60rRlrBplWmKo6kHeUIZQfidbXx55kvMT3WO1wXzwSWkP
GD5CkmKTNQR+Jt4RPztR+Et/Y23SxvEDdfJ6I+W67Lqas05eackKphGXAAHImwLx
apvfASIfNr9V0owbAu97RBKm4OuhJsxpnVV3GBothb4Hrbf68j6/Bmt6nsDa1EHO
XV8ic9yvYxKjOiFNf3iFfKMmFEIBOaw+N3KIdAx/LKf2rUQ/Ysp3SZJGZvajUuDx
zxRch6DYRWObzlqUW0LQMkno4KPMjSqQ0AOTbTAOvyI8mOZK3lwZrdYA3+8mzA8L
qWKYXwJBJlaQZO5w4wMxu+AsY0rjzwcqqwFO5oG87fLvMJpQzK1QQQxnu1tRoA6E
VEfzwTV+YmOAoFyR5l+kVxW+/bL0YaCAY9bTEInln24gJOvvDJTm0c5aX6Xs4H2S
EQz7tSgi7ySsUCIo5+5LtclKdq2W8KEj/wjOoQQs9r3pkMWt4Q8kMAA9yREgyR3g
hFrJZlnRr4FMjHvD61u3sWhySHon4evt84unNzMkf4oYmoQKgpb/VCTLqCdEE24r
LCJlv4uQvIeDSVszLVMstIzwYFFe5PgUXhGfqEYyAJVc6odnUIdrBl7nioxw5qJS
OTSObX2yIFu1tS+ZQvM9mo+RaKJA9+E/xsyLtf0JGV/lEqwhxcPUIi/PQX0bjq+Q
HYxaxsmgcADvLOQU6QOz4XKtz/02NpLZLBARMu0hVBzisY3op4m078THyyEWw9WR
KNqb1tQ7WTR7GLGM7FBM/wAeu4/7vcig5EKn/fqQQcEEijAvfoK4l936W8g2Qqa5
XROUYKRgzNAggbdZvE9hSJfDhJ1Sl4Rur0vkJ81CchRIYXcn6w/XzT+buOY+GSZh
SXNI8vVfnlysgogmo0+X8hE9jHI5fuSIzRvSJmm1/LJlziGDMC2pf4GUtHXNByJQ
LyLkW43Avrb05IoHPEF5fN5A1KRLPNrswxy7gRWv1NkBS59HPGdgSaJtuyATrLjc
7dXc0obg5xKyWG//kqwrfiIdzT7BOc/I+hyd52RshpMVXrutii+YiPwH+uXb/5/5
mGUvt6g9SOvhPXLqkeDvehR/TluQ3QL75V2t5MF0PwYdo8gEE1Nv74Ny7HkR7YjN
IuFdXQ1jtFQ61E0AlB2UyShT5XGJUGJXw8iDPno0nilSKR0ZLVhM///vdm4aHDYT
l4qDIg/OfxW4qhm/X5G8Uojn0XSNObQsdzMllomAhaeH+eQFTGVt4j7+2bC5GoIK
SidmXMNng2uQlArxWoGy4f054G7hAqVRbEo9yd7KCiu+6Dfs2LV8pI8F3RHXJV9w
PGNXtc+GzPir9CqtxH7MCwp+/cUEBSrJYwInICIiP9JgRK2r9p73Wo3MAs7fMnMp
Vc0kVRa6Tfy8+22lW2rkYtVAgi+pjF/IEG8SlzQHGwC2NrCi/wSF1UOFMzlpLnLu
eU/M90vkO31KWgMaq2cCXcF0k9akozKjMOKQru9dvmBDaFR9jRfeOUZjI2BugbVN
icsiNShdy/NRY/3LT92MClEFNvebPtKG9mcx6qIC/0tvDZyg74DfZBlnp7a5Wcb2
A5kPobZDAMvsR6CxldBUvlnuXI4whE/7AuPq0Je8Gjhs5SkI7gnkE5X4CsIflJRM
tAbe2w997caaQN9bfzshtjzUAXJVUlDj7+NjqZMghuYKY0vWptlprvnNrC0R/M9n
UQR7hQ1d41njUAjkfnTECptZ/2GZ12oeuQNTmnq5fbidOJ3rYpuGrQ55EpZC7d6T
yxHQ16xZZPZ9ZqVXo7yyUshcr9aCM5WvtfnszbFkI2PxqHC6Y1WJrsVhdYNivcxf
TdLSSl9+LY0mOy1OKD5guIQHNxr8gPd59PlWggAFA6rn62KtrOwziaR+gpEg/4VA
cGrsu0zVucAcwpksrZ3hYG8VUq18gfCQLebPgZx94FtTK1Pf8Ot5FcanLaHXZ1sd
dBZBKHC8mLK1gDpeR5aDRDBqLjggUQBTFmgZP4Kd9ueJ7+n1xtOLkSD4EGqVjU0k
mHdrgwrWQkXiM49gvsH3fJM3VjYyEKAwA9orphlW0VmTMJ1hOPoT9vEyS8lzuf5M
xrvtYPviZ6AzGJSULMgUP71CaJutAcnVtxvt9c3u0GW6/jvkZEEC2iCfVdOJ0p5c
AM5GvMRQaNTDOd4FlLvp9xZAiyRo7qKXuYSVFBupgEy7Ck2z6h4Tmp9xRDEk32f2
rFGWz2AVas3tVl3oWFOmrdaY7QwUT97uyNFMikQZGrlup68lz9bHS/sWzfYZ77/R
ja0hWe+ue3ZPTo+6XUa/lOD0n721hPK0fOg4OfofXziA5foqI94gQALjeRmqdwWz
yk4Tk900rESu7UTD2Bszgklx3zWgzBpjMIXQ+modQmWQYp9hnhvcgUOWK83++ABd
kMOZEF+9xndIde0/e6TxImXh3QCLJh7GVEt4bD6j7+EI3Fhdj1Hw9ij65vnZzCQr
3uoD90+1Jaw7eVLFLnema64cLt8GfPfQf5omT6M0S6GUBCaS4SdhWKzZSkzLYimS
VD/NK89EK2CCO4PmqMjOvNoiPBwh1lbHQYLt/WXXKNqcCR4NsdVhTLlcVzoDGlPa
/hh97iqH+AzlB95ewcJGfLtYZLz/0+OEfG7Iv9mUFXnazJKGbuYpTBlL1yTluWp0
GZlB31EYo/WxY4CtmXwetyyfGvglEa76wd84W2x1mPElZtkdmJ4DB5UPAKy4MJJJ
pT5ffUsxRcR0PZSevdwzcKwszyKOP4CMyUfKtFcWMEnho8Zog2ySOjbn+Q4F+5+J
IW1sShsYu4EyegvA1Pd0x4hpsTk+pm+qmWtZTSZwLUy0cbZswVLwZcRLlawVZlGc
dWWhXH94MI/s4+y59THFS7lk9kJVRMsUZ5Yjtg+ApHn7DaWhjImA05PTrCHx7BUG
PzjkIJccEQLW6vDWvoiV7O7asCjV9TlFmpYxykICEo/JtvP9NMPPEPtsDQ3OXCHG
UbkSDCTmBqlDPTFnOvxszvVPZjlupH814zdD1HH6+Mi6EMm/BAcOIiXTZTco31g6
lCam3Wh1IJHlXMV11FvWht2CkEL+iJIesOli+/9t8F5Z72uLMRWpomoZCIF4q3gW
DSOD5fNbKPlaZwBqxQA7j46vRm66E9qH9nctCFAlVWxhq+UCHuwoQjKpGDOjp37K
pnRJFzGIm7UO9rHeJVSR6pf/fPJ8fuEOJ09k9PPl/p0NtAufaMKFzsjQy1+5vX7R
Hwj3ctfLuuDwAYywNqvx6zRDmt2yJvUhhnAFroeUUYfVoHMRsT3Q9mrOQ+7xNPjY
EZ6XFFjlUAgxiUjfjH5QmZIdCtb8AQwgCJEwIEO9JWVsgZcFucTQswcaRrqyCe2V
BDsfg+DyjexW4y+Qmn05fne/jMxbP8e9WiLkGrfyt2TugdPtbC3Llrgd7krWFMd9
p3UQcFmFiACe+QyUsjC1VmCsvGIfdGKV2DKp65KeHl0tMvNdPj+F3aWiPx54DR9e
0LK63hL8/USgRoIfuHT/XWH6THi8JDcgzPB+/2IbC7s1/KIpRS6ABrgA+t045unM
nfU2dn9EoI97+ZPbDaQkhYE+uT79nK3cknAACed/novtQ/s4DfKxx4msk7Y0IZpX
YIZrFbKeTH+RZxkVcWFLs7qiSIBZWpXEFrdMfX8DXkVa/Rp8NL/3r9oXIMkOrZg2
DgwpYADyOMklGpaQ8PHDu5EtieTzs2EbMV5Rn0SowM8NinjpFBryWD04DB4KxDtQ
AfoamB99iGtVTx09ts9tGIwQjfYG7pame8GggbbrKej3NKl+U2B3Q8VW0ylYRIPw
AypNuMx9H5c1qTJvdH5Wzt/Dz09IdQuoEtu0bKAlqKxB7e4NZKv0YAanrz5uu8ov
qCDgSk/RWUNtrS5K3jEDtWHGxxvZYC4i6+LLpSe0kZMPRkv01cRBB47gKL8za3ET
eEe34+bY7lxnrUwAvbOYmnuVs5lzxzZwdCAnCdDmGq6/SBBqCdtFk73UzA6hZBD8
jU/cmHoAkjDcxrRPoGZyYXDQJnm/G5SwcG6+3AEw2QH2kjiBnXy0ILNyf7d13aVT
ZQM2Oywc+tPz8iKkd9Xowfu5C1wNdVCpLJFvO8QSzElo15J5QFCyUV/2GyNHzF23
Bbr1M6uSyCuzzaCcbTOuoQh3JQ7YGh3x9yOG4x30OG0FjnCyyiSV/YTllwjnys9V
VnqDkxiQKR1w4C+B6dP9VU5epJR0ASFT5oLaHG89ZGeRNG4jSALCjrjCDs8NvWJ/
bvCC6EMRrWxfmpwwZNIy78jWjgmDY+865mHwfc28Kr9qvEiHzWBy3q6BAloqIRXS
btWz0MsGk/cQVg87enS8y2qUqmUSmX0VMA7C/TZ5LNP2EJvbz6XHx4lTlCnr6XA/
D2ER82WJaQUHP8h3n7fK0euCieHa4q3p3JjrQeDFBC+bHkPHeQ53qb3vLen8UlXR
Ve2rLAnz/RrP7GvFsGBBghxGJp3p+33CnTWilAZ+jHEeZTgS1LWqyedfdJUGsZH8
IEza38FZRdWnRLH9KMF6yddbkdBN0DeuIXp1a4UATNriWYWSOG4j0nBhs7oNvLwb
1izZwcvNCcDr9N/f4zVX2hJ1ZHUOhF024L9hFdlpyGyd/Yj+8Ue5bYOSa6l7SDLh
Uytsw+qnOLSq5pg1tsaPkJdWyeWoHBMTeGOe0Q67uJo+NkjfnW1aAn3GDhZT79bc
WXN/rWFPZ0fzjOlPI+ZndTxpdNLUbQ5bvzNRdk1muHn1nNCVUe9OtNAK4E2KOK7c
t3DQJ178vyvV4NGmYeR49t1OGUpRiO39c17miRDrjY8YQg6g7DnlwGK/hMCcdGIW
Rd4T3lexO0OIIsN/IelHA4pm6HILesYr8yKZXqpvOcGhwy82EBkIzEwb1gHpeoi4
OuRp1pazTCwciW+lU++p/kcoYpqxP1CIw8j19ddanUmmL8wYne5mlH78I5hkYRxX
hSFLHDtVi1OBglNxg6pmwxP5wMW29b0PLI+DVf+Bv6K4xEmMs9Y+q1JCWWC+tS22
sW/82k9roRO9O6ZupVWBHBHFlwVd+bnzndDvYEslR3Ocl76l5NhKfyAPADbQKOiH
8oN0aALj75ccapP6qpiCzV/msvuz0qvPsjHzG/eAwLxI1ejWT8ZwiKbYZG+hdzMh
itRpEiBski8fAxigARUGGY3Cv8ZvLY8mD5I5vCF5egkpZlfb3Eu+W6mNBRTmTI1P
o9Zlg8GvKQSlMT4fBNoqzhzkGZPuJhI/5D7M3gkvP7463tHBJdV1YEFE8DXeoDFv
DoTQAE6rZ6wXMUrVjxs0mhaIlU6F6I27fXb+iQSsv9K4BJiVS1rsVPTlcJoFfrCW
yWT0A5QyzbRe154Eg+M9dqIIL6TXP65WfqU6x/MwQWG1hV3VJkHeszE80SD629Qa
MTKs8cRuNZjDXzlXBj7lrWnbi9Ve5H48wmTuNWiYxN7+QvPOUmfRpZoPaUUJarWa
zRxX5B9YS7Uc4BuAmMq5ywZRU4UZTvlgHuS9eCDJyfrOw45BlVw2y2Ixzn4nGxrS
K9vdcSQIwK0mQCGomhoA8dAaENHS9JvMQ4l7OA6VUus7UabxsrloORll0YIlUju5
6frLmXUjVo45HsLwTENsvqTu5sclooqPjdcxt+zOh2zhDGrxoEj3kygfslwZt+ZA
9gmvazBTJA5NtQSQZJWL3eMn5eDsdKtmEiQ7w3lStMky07thR/xO9WKF/TQ25Pmq
t1Fl/jznTA8kuWHglgCNpFM2Oh8g+oFAEdGi7F1aKatDJbaKTAtZNeaw6P//QbqL
w9TGbZvFIBo1orqyNMVTxOcFRe8ilkvRBbmVwNc13216y/FWVsGFPa60wl9wmbCj
QhGnLp3Ou7r0IzHYccRGRXWFaVnlZiPKfp/aSCwUxHj0BCEm443FFyllf3GbzEtd
g9VSr1wmEFODFqm0w8TNPppnGGI6K3DAlmKSsAv0keByEIgpfkmRG0J4Bw9j6NqJ
ANTl52UsY0yPE5n7bAY1LmNZJXZT4HD+J14vL1erabGapZaplYzwtCvuHiAxYYqz
jfoocb3/4tBxNZlVwROoVSrszqYLfAHRiUUz7QAifJOQrRRcfCeD8uRd2yiZ97L3
LpYxSzxNl9ybjoX4zXZBG3JavrUD2Td1VVBSISkvjcvzgoJt04glXtsqMFfs1y6h
0QKUh2LYDN4luc9Tuov7dmDAwOJVcJ9BKH5Vgjn4+2qy9CS1xJdP4kqyd27kUhxz
RYGGfw2DE6C7zmidxso7RTzX/Z/X0J6iUnUlr5DSY61JXFQO7zy9QakdbnDkXA5t
mUkSLxWgvTxQMldY1BZliMVsBhk0PvQIayBFvIrtE/XV3wQYoRJtjZR7w104Z1wS
48WsM4Og6lRhTP5/+b4vV47E7zkU7beucAuK1/11tCwRj34qJSel4VRLSLKEItPk
kY6kzPOJRB3zpzTFOpAb/qqqgdioqZdWchSYeUfjx1Jhc4jLihuMiRs/xA09hWpt
tGp7EkBMNAPQVdYJZnv9y8vyXkDV3QNBAwKnIXMerH7hRfcxq/r1Jn5Lr+bbs8g8
DndQOslOKCqJJVn6BGHHS4ClDhtlxPsS/nGW8s1as7uPN80ZEg+8923AYWws07BB
PuYDZIlLZrNAss4OTwA2J7d5ZADG3ahq8ZTVX0Qgu9sDAMRMtwcFuPKbhmH4Gd0H
eMK+1iCQJk5eHJhDRHhExwaek871LfKFsluVet5AyrKQjAN8CwwgKvnCGL/G1+pz
P8I18GaNZicjtb4yz6c7HbNl67vPJ97CTCkStIQuAMyS6VfYEbpVgtjR05zeSOjY
f/JZBWHPvV4RozyUAY871ypKHxIdCKptTGegc3G0DnMwDhe8ZYfM2ms/YDZ5/dSA
SdiQoiN+OlkebE+ruX/JcJxg2io3qtDqPGKvU/v5MNsfrPCl6DGdFaim78cC1Cb1
kMYeZD7FKk0ed8wnIsSvfGCmGiEf8bkNNNhmvtQJ+eV9XcBWFZznHqvT4GHiRn4I
y03PLFTMwu2371Qz1y7A/Pjd1tt/aGcuS0CCkq5ve0PE7PhNT7BJFBb6vUYUv0IT
ZZakDXPeNZwnKuFuxCY4xSPl+BmhGBxTHevZmKi5gGBoESdk9VatFiOZv4s9s3Fq
N0HoaNlzTPGOI+abJ/9tkFFZ0o6ClVLIQ5R5N7wfAo0gv99IUpkdGTCQsHnvvkec
0NnN7ti3Z5Hbvzs2R3yHQ+zyf0Oq2WQ8prNFTEcOHHhdq09/snXeADoWLTRN6H1u
3kOA03XTZWe08xQJP2Kp/M216iRk3bGu3+BTECzA8eyKn+wHhZNxUqrRoYX1GZHS
bUZUX1N0OTXmIdxgpUZ7MOvJ/LKp4ZxMygytJ7cqx/wkr02gZHpCLazMxLHauhzc
S7Kx/KRc4bR09qwXHWzCgHTISZlG1iIRD5qbdTZtvjk1IKcQfw94qolsihT4Qm2U
vcffqfU/FwJiErRktYjMmC3pcFrEBL/gu/9SFWpt5i+MY8G8Z/8tNPlUHGfnT/C4
GBn8Dx6Fh+YIsSx/lYHyoEk+ii6q6xJYxOeg2golnlLf0BDip8U/aRB2AB6IJWZK
2fA9BTK1QRTXV1yV7pkpg3C7/7Ybw/5WlUBml58/wMlf19UAV6JeU834xn4NVNud
4Dcrf9jOium7i0TPmbzpKTUJSpEu0rNzjULCwwTz57VJUvdiVDw1W5xrPEjEF0Gu
QWaudFThN+lkGQ01E/Ddt0h3sAXNx+9JHn0j1PbT1ymR/QDSb1bWFGBHNiu2oz2h
ZkRSKUx1u9fXWMjHoLthPrNNIVj4icmkvE1023EUK634apoEsyLqCWgwOQJpY/r/
AYwFdJP5eW98wiuxFJ4lrCZ3XS16TapYyt8gPT2tbqdU/IcNXagcNRBg3YJPz0xm
EJeWgTlNsp97sAavFWcQb+PRUVq/yYZ7U6XGODdGJV/e0ygrXQPDZMKpUWrfvpSV
JAaDAJo82yNVuMQbQD0Wl3nak5hieaa88UaoTBcoj3h0jWRZ+9GjSspJKdIkg/mI
Atz8cHpt3C45T13iYBdZEI3VPHOXETgZ9tI7vM3YUK+RGRTbA4mrZ3q2A9vOWDH1
0A4YJLBfsRf+8RHU1X8lw8KwjYz1jPxz4J/OfUrH2+GN/9n0SjQYQWaa6HnrW3jL
XXoq6u6PoSwQc9iqBkHaHiVH3fAmj/gnG0bxotU/+IljgzJeUgzXaXQdqSqXM/AZ
ye2RCDBH2JXdz59Xj22t9HHUYeI6FHDT3NWyczsa908QzgZGS61R6c6ohc1GZkVN
WwC1cep4p1b7/NkOkU0hODlWBXMRkzgTuEyUOBR81++cmJ7wE4gl7JkOXwSwD6S3
h0Hkyqe2tN5A5e5Evmw+dtgSaKnCmaD28+q8BgxFRSjACi9Sp+XKFiYZxRv4l/QC
nzgHpDmhsufFhw4GdcIb2O9OCrZSSZuuN3yiFXnOXi2DyuDfuu1oWV9+6zYbKfRl
zhczktZqMeCLZRJiFD3FN+r3mi++geCpn/syL9RqWKxBdEjglHzZtl9qPnX5eG4x
kvr3pM655zVIezpjpCGw6RdfqQDOv3GI466eVKjSCdz2RbqrMQSLlHeTlzna4HI/
mJ5Die0nPajHsUExkNhGybYfKey3gexfy0lHIwzrZC6mBE7poPwy3AA3j+YttK6t
oPbjco7AUm94T3Iw0epCicCM9oC1bnaBpmjo0+AiDO79OJEFNXs6dqOj/Kk8DW0Y
dEw/ZP/HefS5U2ZELv5+4+qKzLNzHdS+cN/MiQ5rUeYJSnQ6uYxwuDvVUJ9NAzdn
yOsF6a+GTSkhXGGNesECE5aqCplpoIPEbmFc1rlreeN3cng1jBKMTHscBYz3YZqN
peuWQ+oj089K04W6v02bjvUArymq7Bjq24lZ2AqlD5pl9DnAuqvD804yop1Q3ajK
dFi/TK3v/GyKerkPvIeF1Wxj70TgvyxIaMNEIO4h/Ie7kXvTq43gM1bic70tHfbl
BkMHAcoVn/kYMR5qvRRApGWwkv9Ax7p1hah0PEDOnWpBI4ZibdACGQ/foO9x5sYZ
u5d1plkbmu+2+leenTvObm8bzoKGUYBAjw689Fa33GAtl3woV20JMTnm7QiNHjwB
OMOtZfV/8yHha4NE4UGC5tmOYIzafNAT42b60GhsGI1t+x98t1r/ggYC6vofTx3N
d8wqG8m4BQt9zSlLPoCC/xqHq+7/vdidHb0oA/RX0lH+HaEalIW8zZ8GboBBS4gR
wGsW5CbHc7zDCRZAABijtFd8C7rJQt3vS7rh07JHtwZAZzSR7/xtSI9lwIA2RRdp
rlssEb9frXqNkURGsAyJMMrZSNArzWZ3nVHc7cmQ1MkN79ECE2TtxskUtdVO+P+V
VCDYNAA27SL87d43Alzdb4B8xrkRo1VaP4s3yuY4UNCKi0Rc03jo+pbLcTIaUvyn
p0ODkt3o7tbxRPOaAXd9fLF4O+X6mDlsH1AWaMwr7lJ/oomAyxABq+lMrkn1y/70
Xx+feBeivpbrJezqNlC7PU8EtvYPv89Fv2YX8SeX6R6nAm58QIcCn1gPJYOUrhBM
BztOogYSV6nbeiy3lOZzvGjVf8kgLE1lQbLzesqyCSBLceui9yKmercSQovvG7sd
ZaiEOSC5EATWYBTrR/7xXdsD6XKkY7/bvmy2NsdJQd9R/a/8qwm8sHmo7Y1XKGbq
A9BpaLMQRl0f3SCbLu/s49Vt9jD0vP4tm1M8fFyyxW7ytTfVtXJ5GEmIh1/LNBPR
U8MAwcDfZsgEuHQUhAW+KyhTnekGFJ8KN3pjgaq2yiKx4nFNLx1UeCQlyeFYwEne
xctRha7wV3x3LNYkeCuLvML3fzwApDvobiUib23APl4ZDdYQndmi0rLwCBu/gCSH
Arbx7xvOIMVGrmx/nvK9g2CUBhIoR8eMhnJwe1dEBWXZMQtHrEqErATNRcXweuEH
x96Aq0a4un51GGiLAv7c6PblySthEMcwfQMSdzd9ccoFP3KUWYJ/d6R8PCfNBAi/
opdQK8+wmyvIqTbFXFAGJP04rw4LOxI9D8zp2iH2jrXXx/pa0qvtRe8XnL/eDO0C
DMFHWl6l8g+KG4GGwQnLggAW6lRMoRt2H85mJicqmnBUZES8mFQGYOyF2WnUZ3dn
FwSKvcRtG5Leq4VpaiJcks2dNDzGVBWX2eBbhF3ZESWUJ2KNUr5koffG/1deKnJc
H+EPQBje5lvZQ09lSDCFRG0TIj4LZ/B3kouxn5FFeCl9z/QOgqzODXCgjOjq9KCv
KvXbJbIMg4nRRu/Lcjb8jMUR7SiVmS0wjkWcBAhjor3Lk2+pHiaip1F/0hIj7q6p
Cig9g6ILC4yzDx5VNeZ2LOv4UhAxOaAt6UQQJQAuZAr8kbRO2R+vRuc1qOEJLrH0
x68C4U4vGgGUpASOXe20mnhrmk8iaFoYWJSUUK1NQV7bgYdQW5AZmbUcWxc/bhkr
XXY5Xd1ZF6I02H/PYBqcJEszYxY2lKG1OY+9Lh4ocW++UvEDBTNr7XSH9iBAIUa2
etdKKZuQ7B8HsrXWG3LS3rEkTo1HzEkoFdvk2xEKEniDRiLoYTVDC9j/qzgc51FJ
rMfH0MU7F2I3N39NCeor0Z0NXcImOJoqg9FFueSDTGZakFbNDEx4Ex2D+T3K+KDt
hP4HhcHnWtCIqBwTd/AHVqaUOMYzz9KjWlm/A7mgpED4VnJaDH/7rzL3So4hs2Sz
rgTsboIlohm+g9xeTLyFsoeASwH1niorskYjx63ixdTOPCiv8GPQkwAwHy/y26b1
yXRgHfOEsz8mQ7kx5mD7qwKRqn3jqIZyFhV3O2jC+qf8Bptav8HJCpWraTj+I2uK
Mz10qqpkwQvlqID7khYmbtdiee0u30pnXNHDv4C2KRbDRu3Ur2awHFKz6helKQBW
C2sLLhL6iT7yNad6EJQQLmt8I/YJyPg2S8cuR0SLlEyT4HhQ7YOIcQnZvQ2yW4Qv
ra5SMxX26kCf/N+84qzHoFUBezk/MBv9u2XYzNKvRIGwNabJ9og0RSvHpqzoGpBb
/6HbI20IHbVJTri9Ugh0xO/C21roce3LWEoC2Bm9ANrt3Qj8NQSyqKS372dZRy0E
SuXlgKn1D9sCuPJd3qHSVJri2KekSIp0f2a/QV48LBSc4yfyX6WW1CuAqQzVX2Rz
YX/tMoqN+MG3PT6N1xisXcU+X9AOzGKBPn1pfj7nIaO2KXEouCVvbEepNIKIX4Y/
FnlOuXRHbAk6gwLejsffY4X4FX9OUu543eS24aQZn6V+dHREnj4aZHhk/ayn9U8m
6lFZFbVJI0GtJMF1kvMrKcxZwjp5nNlPHevMK3JuS3Z6xx3sxL/O62jkBKESlRsl
O8wZciuZH8cyhQHQdxtG/SoQV7Ei0rIqaTD2EGyqrAV17QpCfedMtpWKhZJbjdBP
XJJWS+wIJDk8l0WWKeQR9K26b0RKAARyFCWbbS3LwHiozj6sbGLBoQ1+rmLyzJWy
iAXiRM0dsMTzETCSI2HECJlUuzrkUtF4WbWLcf0X4xKTmS9ZcikZhCN+D1UyKu6R
ijkNibRW34TtAc/oC6gdVqWcW20ym7qL/EWf41NYZRomUAgr/XSmyE8NKfLtqv89
3lMCud+ibnREjvBCm60TLz9PSvFizEkJ1iaLtfg4CTY+Gu+vwPgjxZepPy1/dZ2d
/Byn7Uq3wUnDDVx1Y5wDbhAWriIMopJIHREicd1WLfsRqT7Jps6730oERuZQTN8f
MFIN37at7BaYPVUc+ddBtLfjjnodfvPFGuWiPgI6JJ3VAK7i6dBxkTx4tumKXjHm
00T+9FEKi9XeHAwyKqo2pX/8RFHUIPNx5A2oaXrb/a20Q0NcqD3c3vXcy0qJBUCp
HcboWemktsUGWNT1bVw1PrA/pWA3QwlA8DfDO97ZledVXW7jTlLT+1VN05Y+NHSl
PB//7aSgujYnDO8JMKAHhTgjjcDSUoXT5Z8GNDVWfFgluAiVHMM6ypcGHUbXO5Xr
QK9+VNY01UCtFSgTap4pUGXOsPK7Nf/4nY9f9NKFDWxk2j65srpl+7YKKYkXWGkK
dzw5Lcx97tLQtPdQUcjRGxHkTy6aCd+01GlL4HWrrJTH6TSwbEDLtisJoaNP9H0b
VWZZgDkMNCluxIjTu8bccft+Y9Qr3/Tuk5nytsiTalwf0cjkXw6J/VFq+dKz9hOd
kfL3Kh2ISsjlOYf+ptxUwkQOrZjyjuFXkyLFA5SdbbyF2y/9mAkQlS3IsrvE/PiK
6Pg8ehQnbsHogrUSPcrFZ/WlcBgdtcsN1QyBqp96sIV2AUPR9iF/4h+3RqdhSP67
kW0CArlXl2q7nGcrsGoAfv3bCH8i43CPSziJ3POq0LQSq3+j5TJDnS2N/BZFfPdn
uI1UyRZgO5cuWMyY2ZjnvvQrg9nkGvrVhDQZDaU+klIqJ0t04+nhDU0j4tGUxI4C
x/5HkimPf87y8mNCMkqJvILmd9DVe0nASCH1uaYwdD2SfLAP0N9emGWPVsdR7gI4
yMzCIWhtCl3P03/qgAlWT/5/i04Rn2EdEjjeS8VZUBMQN1mWplVsT6NzeFFf+Des
SONeSV7VVNN6Kvskx+Y2tsuj07mndQTG6iNT7sMyV15WXnuxLhZjwnT30RY5rjAB
0787w0vPPYbb77OjxEOiw4BNdT0lG6PUMSMnSAK5Obj8+u20kJROdi7QPxtTxG5b
ZomCdXwNJVG9cIk0wEghmEdWo85vN1ejqCoL/vLulMSYHrHVwJPAzGsqG+EgxzzK
8Wy4Cr0VM6nvhRXjw3KfsNoHQzDYkRwj7ym7GoLJDhensUI4mtIGbAk0Dh5Q8hGR
jQpLKM7jEnuKoZtm7Vx7gD4vmnUui25GNv89Iml5JJWGqHc0hikI1dunIwz49UO0
/fBwHn7zLzENUnBe6PKoETrDpnIC8/NF1M7T7Z9Tf3462jRQGFzH/ryPgrBPqpzS
gcLHgxqvEgOB2VH1y4Ga1Zmgo9JCZBAb0529EMt3Vu3DVURBRcPzeWeHCflZGc1G
sjCJ87DNmhxe5XicWz2HuJGff4bwgbbi+k+VMNgnReDRUPet3BQpY/bLOCptnUu0
tNz+SPN0USU1oeCzomjr3qtU64/7VWv3VqRbBbJr/snnrLKj/einbpKXW4N+O5m4
rZ298/jUmS14RqoMLUHl78eNAhgguzOQd0q2/uMUxEM2MoHxoRgfLEJoLw8lNuG0
Q7Ht+yPOIEp+T1lSnonU3FRPLT8HD7wOJwu62m2L9sKEPN1H5K5xOLg4LwDno9GC
3FxGyim4uqzW0pjluZBzQ7L84FdA/3dDoVFkFG79KsKp1YNOIrrJACb8bUj4/l4g
EsHuq1SMpL0lQhoCfiVNxU8GtCkPVeA9sTnr2nrYP9KvNQO/PRJTsqocsZ8Ie+IY
T6jgLcoJUDtUzQ0WEZXvH8yaee9Dzxbn2SpjjFrkgucHB5t0ra5n6/fWnzRgiwRQ
lp1t77ACL5L1Z/BIsnqBBUXAO06a9OzhmfC8tgU5vulFDb+c4b6TmLAzNGLmrjrR
yzsiCwSRm2qkdzrC2XRkQ+CAugKkiZfCWb7PbMhzcvb/4WkzxxFu/8vvcHv3kW6P
NZDi+NQFljvZt+q4Y6kiH4y9/jsWyziCp3Y5tGyN06FAP03KSbfOHYuLs+RZuKDl
jx78U7+H9zd+aTeZKmjHvquOJIU1+k0PG26bulHqq3TwO/5RzrluiEOWPLATFyWD
pqmCnVLu40gMK3aWPomrrfmbRHIdI6ud3AL5b39UTGq2nHycrz3ZD9PxGiP6/Aab
IMjbJK/g9Cgtr5veE0tLotWQnLiiIiU4yjb5e0Wu90Cn83/cDLypDlAIuPJJaOFL
04itoqVSWJeZLf2NdaQ0NTOEAkQWEVM5QgTH9FRpZo1X3BVu09044AgXKpBl8zAU
mIB3Sknle/NwjHOosJ4IP5BfQeohxnG5JL1yXJEKv775Igkz4GiUqCBwHwx4TM4w
RXP4GXr1I/ZGXmiang9mFvnPkilxgklFZdDI70Rbn0wgb0i6KDco9KQ6WASDDKhx
BtlCu6gtE1377bsq7YoDqnfwsDSZ4zcDWv3xEwSwy9mvvwgJSVpNF7QWQavNQu8d
It+Rnsi2sJZ21AdNlABX2pxCHihmMmquO6bUftAaWgZtJPwvKv6quEjK3AYtTWDg
NJgwy7T2iuJ1C3xO0+n6HcZ1HECJipJDVzwsLyr8jhZeUJNz6BHA/W0jY63KlmZd
w/sghwN4RZ2gI6yCJ4fFAOJGkxyTNlpRMwASpKA/bF4Lfjmp6e/M2789GD21Dkxh
+UR2HoQc5YOFsXsC5Rdb6xBxlANrI7FFkQmaH7caVW+p0hvDJ0Ekj1l4iM+2bLs4
bUvKgtHPaL69mPjAlCAKvjifBtkUk8OAl4fLQdJcc+wv5vTNu50EEYqpc9UdLg1L
QQfU+kfiI3HPgpxnh/k7K4b7bmbHFR8Ed/pXLxW5HRtwxyduIrk59SiMRPWPNsbR
uIFiNMBmlTuV7RqLrheBdF3eI2wPCKIsXEnC3+i2u1XJ7HuaSXEZarjQxZxCuA3J
9x3v0/elA7Z1D4336cl2Qze8Amd1596ExJx6fFBZRn7CVp6El7/NtVHK8ms+KWa+
nvsVO8XHcs/TulLQ1iWGUjXgNIeNI18tJxEoJhZcy/YEOFlMXdHhCkIihucLIaq3
f9HReau94bc1pU+Q2wOlk71emwvWe1Vjcbe/LDbO6Jocq60XF5S6Tb8dIIqlLnWe
HnPeAsPAr+3WbXiGwKDAz3R2YLWftAzps+IciccpIWthpOe1BwVaSKZAa7df9GLW
PFuLNgH0mA9NuCDMGYy+ktHCC3pLgLmMZfwsOf0Lb/NaceoDF7+ajdOoEt72M9iK
CmgSBqAp4Zo/rOSBFNZfgG+MwC7cQNMVnWNrvY+j8YSifbR2EVVznxrsdr2xz/k7
DF95CulpZLh6X6PY1IX2OSBAXcKRICNyBbt+iho3UDUVKcGsa2Re/3My2xZNXLnj
EYWm+9nER/3OPRHg2oZmpOYwLwu4eKwSIRs34tEVvZTCM+/WyZcpCgTcszI9fPbO
Yz4W7DCeKk5kTCXunxRRyt24rXqVjhCidNN6ank42rIHkn6v4J451akMGPbgWkNu
zkOJoMnfMhL0ZqGdF0fs7RQ+O/T0F/BQwpNSWWEbwRbqtcWdl2VQtZ9+UEEMAp9+
PMxQfXchDHQC1I6Jp0ILZxYGafrxSLG19YQcpaPem8qBM1XS2tBI3I0NkrzqyEIs
mhrA6jxl8X9gFufN/3jhUbwBJc35r2Myexk6OyUkFF7c0EwCjzVthLGPlsnaEhwq
hYbvBN8gwHOCwpNizU4ulnOyr08LuvSZb7eQHs2TAbggNUuE7zDl/gMSgb6sE0vH
OYjNrkICxnT+gd/UAU3eLkQYRks8G3FeMPu6LupC4HXH35xoEIo4K2SIvbEm16lJ
tPzwVNRdC9TuySpRZ2q9Ws4006BhjhV4rIWmJywdoLbbnslgs9vKz2AOM+XSwr8U
irwkVftrK+Waqz1Fkm6FoF4ZDzAlXMza34ANkbFl2VFJ1EuNj2Kdt2PiXvP9lXiG
dTkj/2cJYW6IJqGqx/eFZHtO/oaIgCqe1XPOIwHYksZRfwb8PfGT9NNoeJZwIBPs
osVx/BF1QFyDRUk9aPCu5JXNdd+2rYg/6DMSk9Enspvy7nAA9nhcg7pmchxodDoV
ZyC4WiZQG4K6zl3l7t0YJ/hzvgACph4sUaCdm5J2UkMRw+7RTV39BdXRcaYCed0g
EwLx8QPbME8KHGxZtnQnV0tbNp5NztBpRRAHeTpl65dxHtIl//VauxxriT/qdb6R
7fcAUBjN3jCl39o8EcuzUBPWeiPogNOoUSlbx9ji55jrDv2YAlCpWzNthzfZ8QB8
i0ZtKIx+ealhm8QHanQUgW/CS4GeUb+kS0whTeUqzgkJ4uPWcfgESRbedqSZIK/k
+wgZW9W7GQplPPF5ao8zSSsBLjCfXA3Vu8Hp9lCfXPySpqCYMSejxaMzqtTWvFEc
MFlyBFJlfc20sCTA9GAONYnLS3vMubbPwOOFfUq07jQqwswi5xguisav/8N4uHcB
nkOEJW3u5wX3y+kf8+jm+FJGqHLvLP8KDxy8w4BpdWYPYx+PkFe34R8RISvrnzAU
n5b6lHJe2cHKWN7D3Oai5NeWxW3YbHhAWDBR+oMmDSuRPfrloIZTon1Alic1Khvz
E3+ywYUgrsNoGCqyHtdy0wzE1+7Z5kJ7BJ56mZ1REptFzn6VMiT8IhgIf6IIjWr8
bk33TQPcf4hkZpTT1wSPgsAVkWYLhHo30uUyft75C+Qv9pXWwsFVq9b6QmHdY9US
Ro1mJ8sIrrZDNIyoJgjPSyVOIK0AJiXdBCmx0DD79oUOJOMONmv6AWSujrbkTvbh
IY12gYURjoqy7kgxrWyigzgdhCRZwIBZiliQiGp7HuPyumCjhrqg+Apth++tfUIT
wkpD7yys0F9drImpPa2fnm5dRnjZgs5RaurC2RlXg6S2sPQO/R9JgnYeVxdroFTq
DlyIHICNBcVcFILTm8BuKcDzRq0m0fjhy7f1n9ZEFU3xbNUrroonVN2Ap8V/EqA4
cFcEd17RyK6zFdL+/7yzenZXa+6RvNFPqVFWacE/2yNOH62oipibIbS3Y8VbGyYQ
VO52+vHxH6tpf65evejJriqhnBI8oGYNxUeVuqyOUUC0cFeATCWK6CQ1HkF43+1I
/RtuZlzc2iQMxTpjWKkP+FfWkK5/0GDT0IMCEnKH1sxNSPDClfOD/6qtXtxLY7eZ
BRcazzqUbMO/PbrMCNqtu3lzjhuG4zAbEyWsToswHYDag8tr97aHJvq9llajscUA
+6LCYfxRjfqWjhw6tdfbc60IlG3rskmSXlsoCR9WlVAOXIhN1CXFLbdz0DoqbHva
Gwlm1JWK4iFsFASToJQISGN+7MBLYim9zaB2QRpIbxMe8tP541N6jgOKTOE0xrXN
ib8DmWRXaglG4QpV5BWYyo/f71qZeTiS0ewdONCnAUpHGvkCJ70sA7vRm8jVaSyT
XfiA76ljqDXFgT1VxeIANzuF05ar1ARbJP3OQ2siAQmdPSK8r0FU54vV4U50AOGC
hqPfgiyc9748ngg5yokT/a2FMPgPt1J9yzla2XG7TVs/XI8nGo8qs3tg17Y3mBMW
ksoyRFk8GfzapEjCcndBMG7pSPsRPrw3QEmSS7YPYcLsEeM2sf8haN8r0Xn2DjVf
CIw8cqiyJ+Uj13tSQEUOBj/L7Z5qtQ5UNMlXRFmyr25/PH1O8gs2tEE/bSvlFtFy
5YXYRpvAvg4SnCAprMuX553iMJv2W8uD5U0cnEg/U0QWHR069YPQ548qLI9pw+tU
DjzM9VCHHN0WIoKEUGfrzVOw7a0qJxRdmStRcQxACEuEwMXWkHi758GjBNY+suVG
G5+XHR2JVVdyNs/kzSULzc5oGyuizaTaXlfj4qT0h7A1QpVfUoA42uCKXMMOlPsP
/oVU3ptE/FBvtGzDLdPkOPsgApikazr0xxFK/Nj3LMpXBfgr4MhG2CO2X23RvZG5
gz3i3EqVOnDMbTmYHL8OXSWwYx/Lhp97gtgivQeZDF49TrJKrMsubOXq8QYKOyuW
6d+5mUEEVgLPWJqR8gEKyvtp258Peb33tCFC9qTukIZJD3CKJHGM7YUltjNimhg6
KGCgjzkWYpALKiKVBgAQ6mp5amHznxqjl8oJi7OeB+GPCTNIlCZIwaQ6lGKSPQ/s
BmZpE0IeRgDD0kRQuHeVbLFhhJcZ5onHqj2BkeX1Grj+YwzT50ZsCeen+TELfLmb
WG8deXFNnJbxEGIjng92VQ+hoplgLO89UH7y6YefgHb6gfvCQLWkaXPU44RKEoeu
TtHliEXxhuN0imXHC8m0lgOMSauO+gVHxOqp2HYPCCShRc0kYCn74A9g1GoAkpMj
PfmwB3FPUIxtGHsN9af5wUlBDS+k5xGcdNa2NCk0OeazKyq+gzBnlQGMDD6K0U6r
ZEENFCXhtxwl8EWLtIz6TrdNOqwHAZVfQV2EV8MKw4n9jFN+OXUKLScA6VQjuS4Y
hz9mRujEHUa4OQm96M+Z9EjQIlEx6bHDfUmSNTIGYDMbeJyMj/6gupyqdVY5UblY
ZOBR2HJtBp43gK/EbbT4jURyyA1zn3H7Px/OtjstsIbA5u6z1mRtbEfqLGw4JP1f
av3jTnnl/aHIp2oNfBwtzgl8mN2YS5iQTrM/lJqxhQe9dtEcyfSBQtq1Auahc+M8
85IQmo9/uoSgTbmR6AR8dqdKOgd1iCnlA2EcsvEb24PbFe6fx3ogUFYOBjC/HBv0
TUKApu/XEFgM9WZDdlfalqxMOplrpsYqdx2W0flkUp3Zw5kYBENAFfnX0P9vtR9F
dj7987AgGXY+Mbu+ybIChjmkM5EJH+B7+5nd7SinanBYC/rMyVgRX1nOyMyARJFq
eJ4kj7onXJGEuFALgYNSvtPoMo9jKnAS5pt9qkVkkuwOPTxKAFXrSxF+EonA/3rm
PoAvssrjn/eJrFxgiShyOxgTEbMeR71YcljGZvjLjYpNcqmiTTNk5WGXKIDJZIuh
bVmcJtKqdTiskObCTBw7pxAycAlYqkjviUC1URzPBE8nPIven1fXiUBeZ9aX3AoG
khW/i5wyPaQVE9gRCH3wHCB+QFNJmKtYaPpPopmoIglOOsOSZVHJZiDNOKzZg2AF
7jtDhJQXeqLBdq3mBx5/SZuADma5+qqTtip2vR5ukZiJlx1daT6/R6KPTzJ3SOKo
e15e1NXbaGS8w67UTeS8bSwy2tXrA0jBlxXEoP1W4VjyGUsv+xX2XOgnWHWmRI6X
RAiI2v5vCMQP9a6ORcBbVgt1m71+gMIC3pmjSlLZNCWiOUj2toWIqZD4+WThRLw3
83yW+gq7C6K3JtDHNdTZ4cXVo6qVbwTC/8waJOZ7ZEoq1opFaRgRfDQeUXhpid2b
yjyjXaAOCejXSovVkw1rZElvgMlfyNPbOVp2iujKlUa5fNA3YcqVYnaoC6oBfbUI
EB6SkNpMpJs5CxOcDj/s+mdZe0OVcqpIS1yrj0oOz8SNfwubWH5tjDz48H3GwTW0
2gdqV2620Wam4fEeyyIWYJbcsuzAMd4HBL93mX/gmQZw0sLuvG8/jTeObI9+1The
urLc17zxjT0C6Yd4AaV9bT/2wReZReZvDqk6bfbAy34mU1Tvul8neIQQQOO1aa8E
kWc1wTX8n5itV9kpsRtAOcKYYdPZ2NFRzmrbtMlqjpETXhBLyqUbpufUutlKYaZp
xY5vzQr4b9rwmhoyRrA/32jW8BdtQcsFDM+Vmtz5zzVtCK2YOrazmOd2iYDDtG2m
laemuZh4J0pvqHQKb7ils2wC9RTGwLwiWl8ZTmdXdI74MI3lnnfX7Nj50g1Md361
N9I3EC3704+FcZJERt56PcOikCKNxaiYwa4n0eL2pM5j4exb+nypeNoMMidXEeeY
3dAlMogVv6Z25HOlXuypcbJ4yaTM8lYb3cHWM6yPWWG6QNlFYCzjFWVvETAT7YyG
1U+QL90sMANphkLfHsDQoXmy5OyRVQxjCZ9XT0n94KuTUoHg7Kxad/liy9A3tCvP
qPe4+eNj/ZceFieYttLpfh/+NlvMCGc7Gr3kv4T2KrfMFF7GW0aTInD8Bu8vsoxi
igcthyOnrzZIQpgmF3uLvvqtu4I0tBEh9dgPlyumBQEIkhFZic87BP+2ka06K0k9
6+UqvS6hnfNr54yWXMnV5GUxVzGRy+7DIPZl0sKwj3ZL4u6pTD0j6Spm0t0JOYmU
YCW81DJmyLGuvRU7C2QQ0xlYCF75fCk/cvxf5G17u4gnFPgxT11FtSpeSKjzO9d9
QisKU5Sn7SVGvBlGYQnLzy2lBatwUNbE6xxU3AhJChK1HgSvdyGknt8oin3lUGfY
Lf4yCWmoV9saN+LvZzgSVr/E7oP++sCITWwtmuLerhvFcjtOYnaFOKmuLac+Rb+1
rgHnlCEUbd9kzfAXyKRM+OjdHMeifo5c9rzviPK3h4cZyonNl/Ud5ffjWsg94lDT
Zn35ZPBx04qRMhVDPOL11Z8SNtFvaCKD74/Mowgc9ptJLV2OHzJy/qMuwAKu857a
qWlJ/NZ1NhWVVpmTNyCgEwB5rG6jx7TvtnABYh+piEXvJ4v+GFOfQ26ADLG2jj0K
P9To5mfyWjKj+S5Gqan0AEAObyEdMHitS8Da/ET4pamx2RbttuKEmvHzff/VUBPO
GMemqKppaDq1JVV9UISAy/m2SK++Du6W1pX30jHJIFrqJhRHQIhugQcMb67lHsAV
Fji+JCTfT4GitRuyrSfVDqdPFnlvXU2DlWS6tCk53ZidKTkx+wKry5XhqFB5NtkM
i7YuSuWj6fNyJd0LsXBmuocz2+28fns336UdtR6vHg/bCjMcEMHan2//n/KoJ44T
Sgg+wVvo2f7PJ/2thc3r2Q3Il/JunKYyY6WRUSumKg0jFVRix2sbSGFzlXTqH81E
Lc8NX3vB9Qk25RgrGaWz1aEFqaKocJrdOlQG0phyFIk5g8/UBeylXhAR6ERCSgwX
fpeAa92WTBkRR1hEySeAZHMsPTQ9RUkC+eudRPlPoDYpNQY6F8JYowmo4VTBEX4h
5KMNLdZe9RKfKS6qI6FuX5FE12sBIK32ePRF94PLUZG6acFGDFccLs1VTdooILpd
tjUzP+4CjitKN2DEtrSz9dpO1Hh3T/H7BIJEdqq9wZlJEhbmg8hPOep9BH2XAHY1
bpYzkzzRCkf3yEVKUtM2i7bV1OX83nw7TwD/zHAjsc7Xauzre4uVQ1tw/7hDeJ6b
I8SFHTGlKRvq9fUO4LV9RETZnCjsmXOT93NHuqSmvx80lbaUIjqb1o7JdkTFyUUS
TXsJMh8cqlIb1Lr4KeWIqJL/5mko3bygAlnwwkGhKqvlLIA5O4mYWYmMOQ7yZDC/
uqefJd+mGnZXAXNq1J3BAw9WMguWWCLusghAVSQnR4vUUErRpQqfsmJrPF6ftpvP
6KSCNba1VxF8CJFJWofSZyWFirAaehuCAxPqZ7aMKo3PAx1Aaa84ha5Gn2oUyclQ
7Ct2o3lZlm6bsowg5rRVkkX8wrwmunjt60+uG/Nw3F6sGDK3j6e73vd1e6nol9hj
BWBZnpjzUQrUvc+xXR3nx+975ZH7TVvxC7y17FdffmYaZZWZ7cwKIByvzAzFuKXs
OsPqwnRcwVy+OXnCMB4zEmgKCeA4yFd+eV4rgsE6cLvXJ53gJKfXwxi9XJML2nUF
BE9TQ3aJA0cp+qJa1bgC8LFr0F8DmaqQnC3nX+qOUixYqYabtUjDLTZTWScQMP32
7tAj74kNNBqC4RZTrhuBKfKBaB+db+JSML34RzKhaGJYOsBe1bVVGGtGSH1xMIOr
lLgjS70VmN/7dDT60cnTNLKfroxJKP/JCQEo9f7o1Ds+DZz1nH1tdMvdzDuCMfR3
/WdpLjNZT2U1ngr6LNr0Eewih6oIuJnRSM5Nxj7B59F97/Cq0WFQtHXhb8K+xKRq
aC34zw4me7tglJRB2vhGjuON/XJ7h1k4x3tRbeCEbHPI+8eRkFVRT+VDbzpxSFx0
eTPhYXSb7uESD56gzEZFM33HNV5CogM1zwZRYEOUwzTr4ORjVkhxaUInf/sJbqQ/
Bq8onJj8IDvEmqbeCvRbexYTgyjjfWWAjMEMVA2kulW/5NcAn2WRSQMpamwL1ppB
xCui1vGNHoCIZptuxodlASDk3x/OksarV0p39Yq5OdhwI0M/nCn9mG+dfKtghwgy
SSuLcxwRHO1oYDLR8ElXEJ4TbGOkdzF5+Vg16WN2waYT7S+mZvSVnCAyika1DJNz
2kF1/JwJu9ECocG1dARFkUFGo+FP5KIRW/Ztn6AO5v70o9dNSTsqQ0cdPrctSYkc
NpV4sJSZdG7lY1z8zkVe/S8plwVjX91dYMFClvmyxdEHUgLIFVEVeDVBsTCcCSHG
8daFUWa7qhXVQV64eLOjf5tNvgbkWDS3MAASJzwzi6F0rs/ExhPnGZgD5gwdM90u
YQdfjpWZcrCCPx2BYTs0JOeryAGN8BbTZJOpmfDA5XCm7pQrl8voocegefP195DX
ajCRNl49NjpbZx7Ua1Ox1y3Ot4ADaOxZjeThAmautkUTHhywPRoWZ1ynmAuV3scd
sqoZ5nniJhXD64AkzjfP6Z7r8LiQSOp2W1EbGk+A0VUX+sMD60GCCLLD6P3Kt7S6
3HKQo2Z4wG++/mbmeidydKWxwwJWgBwCS61TeZmJvw0u5u67Ynp3oRNObnchHI/4
h2Ewkvn8zTCf083bsuphjjNxlK96lUKM7Yo/B38I1DShFza0x6KW/wxhEyJsAJ9t
qYNq7L/P99OHKu6tjQDL/Qnk/iDr+CqnhCUO4vfDoOvzMKykvr7QqdMqYmyL4Fev
jD9+04/OY+UDtCIRQ0abN+nA1sHblVxJKLyoyjRQo7TkHBGx8Ct0yS3/IUGgSNrl
vJ+hRlZtNsSQ0refl1Ak6hv+rwXerVgwjH10o5uR2kDZjAOIJWtw65LBdrQCu4fU
Cb0P8OwXwodpMTiYHP4HTA+WG0J+fRWbEBxSFvmFdFoebpSixvnYQWk8OUmKGalF
qVqvLGZq5jqNyn4c4g/ihXkthF0YQVrhfptIAYnQUJLFFUd0QRAvdKXZk6W/Kxv4
zOZV5BGq9kyEHVAZ5XC28yJN4h1MBP8m0XHY71/20Gyvmo/XVszhkyoZq/Q2gWz0
UjUETsNHc1DfmZaqeVMdKYrYPmR+japjC6Zt83WIsnPgDK2Pcc7/nNyplQtx8Qil
ueNzTJ5k632jPoKKPCt6fzFPGyGdnEFPre+2k/9SME4OoOp4V2F7H5JYo40N3u7Y
dYj/GCw4zsbrPWiEqOEL56nTgd0nWZI7i20jyGBBv2JIntNTsOcOZVXYZMhnr4ac
YzTQLdoYe6Ku1EWzWcs1WCXfhqCKCMqONQ15WXNeyJOwtY9Li/Yg2p/+Rpfo73lg
HI9sDvwEnLbo+MyELu2IhvPB8jMivkbJ9OnMLHHeUSEyRLn5i+PD8H+OOmzBfFVe
0EDMWeXIVhi4VbiJBk7y9lipbZMLx7PNF9ngo6L14we7L+XQCmTbR1mLW/o8KlZm
ygJzt80rmw0QgNmcb/HvtkyAP41RaOSKTIstbHAV0ddinPULUk/xpEMuaiZARRTU
yV2Ta7Vjwd0jgpebVH310t7qDyaCR6Ao4chCl5OfbEc0XzFj7rNwf3naqeeisbAL
YmXC0blO0guBK2FYBT5eELRjDdaLTgF6WmUGXPUJWgyr1AkMpQeMGeMcHEo2gS09
K79zrKzTeXM2bmZak44MilrVfKanK8Q+HB32s5DxAi1nroMuZ0x16uCaKsy6mG4n
uaLl+4X1zdcR4OBF1Djw8HmFMITXczUnssDfMr9NH2N0djcSs3n6gb4JfIitFbsg
W4gsIw9MuFOpjrWU1a84UH7TJ6sLlOBgecRY3/c746r5zCsjKfG5l46zrPZkIbsb
j9dA3DB8pYnyHf/QNa/fg6JRHiJtYwbbDq+Lif+4stWVqsiSyK45E6BZ2yBMbUOg
Qwg0bWLBhVIbauW1jQICtldG8Ogxbb29qYVdejUTlr9+F5tK3g7igPR8gA3XLJXj
Yr7Uy+5ouse7+8texpOyKFzfGwb+uzcd6eLbfAbjg7Iezw1FL8PU7jnow9Df4CHj
084/PKJBhjblgl5mNDy+FqBRjnLjfOnx1ZsW5/nOBeWRTNCjbl47W3Gg6hVqIxiS
x+5Sved2Llbw//Otnvl/J0Aw3JHyyv0F1OzKhSMBbwRRxNlHAy4jyqf4jVgrdjEJ
MDyfcIPXBvLCRL62C3j5oDRf4uiyLjS286B6Lzoauqt5aU+43dhBBFf7zWgRGY3n
MtuWTY5RAU5Q83n4vTrSeZ2hQpSYyXQBCNZKZSuN+HWv1Rgm0NsF/w4fhSO8oNoL
2Nq0brS9ZQ6AZEVrfVH7wOM80QDAHRHJm/6+vIiPRO6F5YRMDxDIqj5/EuuuBNE0
WuTllyOimQH2mvuBnlPTAkaybduaJO0ZzAobxI2DMvPswNoXAFo03U4wdUEcY50z
N/tGQf/DFCqq9Vv8pstQaT2jdYUlnzV9L0DW+iAnmta0ct8YpkvUnw8STPaqvZpW
K9+27uzWFIOyeXhJX+oh8rl19xkzJFV8VNtsAmZUjAVcCFFjeYs/mrdy3I9volQM
fEulLyxm7CrbXuXKDlHuW4/pt3HKmG/7/F5zbuP1bfE8Ng+JA0e+FFhzwv+HVY6k
poLdjgZYLNC3XQEHV2bO3iFa2x8tJy8nkvlfyNYjpcBbeRhZfNmpMudFBkE2aK5O
E1NepZPXkr3qptUroBoQcVWd4B2D5Po2uANgb1mKRsmAHbG45nhB+FHv6tsSrThW
+iq9k0c7OImlJFaMZJPQ5xjQ9asyD/t5GxfBRHOjz2QxMtDcHQeKENsMOZlhbi/p
bg8aIrvgRnnFQ5E+4xGCNBBBp0yfzj0vsb0YYty76l7dOolN4u9QkI09XPKe9uNY
geqr0WbzCZO2l/jIPtfsZrFjNlnqtgRgbaZnut3SFeN6K1mFfYh0gWWMlpZVkMx5
iza2HIgkzb0WOdB1CMICjLYf6OsfWQQwbn+GF4vAVNLEJw4dHmuMHbC3gie4kKpu
KSBVOO3l9fnQKE6NhrVfzH7TOyr2A/pPMwbZ3JYmFErajAfAbBhL8704P37eqi4Y
KwIIZ7/+Yi4OSA8B6r/98A6Pz+woaFFW6N+qnmz6m1OyxOIskrleG6MknvPWw9Qd
03GRrSVgdoDcwXZIBfri8OpSazzYnZhh23GsBJ/6UXr3Fzi+YFM2E5ATDn6BOJ/m
fMkfbvYvteszXpS6cDKGPZsnVnX+WTTwjJIBWIiJww9ZdYc3W6zEsgvhs4D7RwK9
lx07QyCcfPXCvw/DkTTQqFuegARBzVaJXNi7hYr41j7nhnfyr9S0ovIISomI/e4f
P7JU8Cn6BHaUS619ov6Z7doH56fe94UE4NuMbiZiEkBQps+DbHtv8jMqanf7+QuQ
mP6UYE5zl6KSnala70/y7g7VfT2bS5DIwmsP/tj93Zv7z7u0q7wyqXFI7AB5p0dx
wjJ/I5HEcvRV2SQLAmEO1OOaB6GiTfRydZfjFidiJyjqcj12FfRpEMcsHtS7tOae
s31ymXaQoStw6XEfVkBfR8ngRYjM/G0HR2GJFbR31dN7sgRwBg1H/6GBa2VB4lqK
6mROBOVzPIiDcNpALb1lzD7zGRpWcBWRknoOULqdZrUY41QvviohDc4/vt86H239
1GsPs7/b9WJaq9mzfwcU/gYzL6Ge3gQqpXOXgaLoMXmBFo1IcZgwomVUjrhX39Xt
u0s6EfGZDxZ/o4fDsFiMQ0C6yIiOoyRDT9P7hmS95jDVGYIxzMw7wF/q5mKkejOg
0709sXzzYDhfe3AEhwQmEu0QEMZs/b9RX9l2nnke+oPqVN4b36Tq7Lq63N7slj3U
ckOa0dS7g6/XmHfpKQjuU9U9h9NuCPjIXbQXatbE1Kvt8yTpskST/lSEFma5pIK+
Mvnv5YsCXctuvXNjL41QYMUeFjDwhsow5fIknp8abGxR3YtQrQB1YjZWMuZ1a7pM
d5m3MAhlNI7uXCQbQCy12bGLqVVskd8oa48sdqcZw2zZQXlDAhrrKvTgvLh2frC1
ElQqVJN43yM1zGzjwMyoo8Tey7t5SqEOL/6A1cC0J8rsShoxSb8Uhvgl2xjUEi0L
4/Xwd/iKAw815xZMtqBlG9Q6/SpUeuKku23Fvy8tAT1EqrGhTCxqtgxnVILnFNc+
F2CxQnix9QUniilvPZxLb8IM8XIdiqAA7Tl2UM9uKoKxvYapeStKgqMjZm8Ez5sl
j7S9yhl9R/FKrGnDdE/XvahN3RxKTOrxdz+Gelt+GxAHLiC6cNNvCMZb05O+dS9H
b0gGW7mXT6mLqKEVR/u1e7FbpXRN6TDUVX+XclwN+rWR/IAasfsMV7D7QB0wsJMp
4TKLlJrRW76bJ8ZB+zZmiLncX/eY7h8QzwVqpwV7fykl2QYPp/+IoIhcaK2mrt2S
3WMemhrNVZi2sXAq58gOGAEAr++bmVHUuHfGkGVwXRgQOYQp/VT0T0LgexgaacIs
HfX25FfnFjFfoH3+/m0JT+QLhv8yf9HHi9i0d8AvfhbuLrzNmSwtsEK2Wj+5gP/N
HVm49XoizAuh5ob1Mbvr/tAzipjqGmB6vAVUzbNJ8oA5Lc6zGlZqPJj4Z3Jtb3yT
06UTcCvekyt5ZnD6rF/v9YQCAAGsIjgTepFCGpLxfJsDayKhs6p6xMjohqYWhkmc
KTnV/q3qnSfB9MTq23E9Xd0hdHMqzw4ORoxa8nu3GYpWENJ/KgvYB4c2rp/kOFaU
p+QyTfRcgM8LtphzcOh9XoVtO2WYbPvcmSK+0NPdpCtGR4IVSo/U17j/5Lf9vzMU
rYpLn06AtgPW4rUBdvlvTjcXw7x4D2k0rU9dUCtx2m5NlurE42dqW17B3mKahxGY
pGb9pFRrqRt7zxVJOyHBxJ5Gq3wjsq2/p/HXSopAMjLUG0QgVCu0/d9OKeSbRIkX
wn+Un0cJBrxWEXy2n1HYL6d5b6IuSZ/F74sFyNDFbGlkoHbNpRBCigSQCj9P7rlI
TYjjiMvW+alVX1gUMsh4eGDqQYL8mBlTMP64GHaPdSFC454xflKGYB3sAge8KSR8
tdPAlHJcOpAPCSX03ig3sQc6B6YhQZoMQ90x0NEA0roFFkaR1BoJTWPMRsvnZIc0
tOfLj7F7uH1p2DR3xfi5Uh4YeFr4YJmm5pH/+5h4r2hmKJvoaNx5oiaAbHEkL1HK
YSmF/DhMQAW9Bb+O6Beslnide9z32ni915XsmeG8BDwbRcsorrUjGEi6KSh0VP5B
U2StbAMLmBDfjvs9yjxGsrvmAtc3Wq9h3JOTk4S3u6AWWiJpRDnM2mLu0+HetQVi
1gXf6sCYXqeKIuJEsijkkOm2ECzaW7q84qt3lU9aXyR1Z0BIqambC5lGk1imQ43e
jDXhwC9ZV8mDpviU3P24kIFJM/yuUx50z/8iSyVSZ6Wknen6jnVMSdlKkkBvlLUb
E2Ba8g7aFWeszFLpWKSrS/7SC99qN/DBb8FIoCV6tyUA5tQaZ1rvdZ6j0Wi7alXc
upF2ttpF5Gran+YeR4Ki7yjch2ML8AS0Uoc36XGCOkcfbLnKUuQDx2yK5CQsnygx
cIRuN6sMVUxYsqamcnVMdS+C6OBrw0cgHociDUeQbJDFTR46N7UrEEcurcw8XVm9
1dZIpEVf5QpZEsVYbNQzD0dOpoX4MAyNLPMHI2SPQpit4P/jcQrMzalnkc/sy/aQ
IkBYz9CT8/HWTjKefpOm432elyEAEKA13XsVdenxnOcVULyhCjmjPpGRVNNWi/Gi
3JaZV6nlaxgCGyFyxtdg6HbOjtH/EBAM8KIPWnkd1eLsbaex0PSSZUj5fWlqGn0D
PJGwoFBg6oEzTFv/wSglCbYnV865jEATW29YRof6wV3pCcUyMM0BfD9WlvW94S90
AYLR8kXQJM0xb++d3X2CUsA+/lLJT/eEP14WqzRSsiynKNg3jxMfCg6UmrD1vF6y
NdCP3pFhg+uzk7f9hL+S4HO5Y5RikMd6BEUW6TVrN6uKNN8ycoMw0f3yYZtSJ/p7
zp3Uuqo1ziF3U9uSs+4OoD31+WwwNaG9jqsm6CNk8G90C/XdIoUaDPAiSRrDq3pn
mO09ILvlw08GYi+Ec11rGKz9JtFOLsxflfS+JiS0IRv9ld+TLlOzvd2eVekz/nmc
2VF/wRkcuNAgx5BdZXtf0/gF4kXz/wLgVPSGbEdF2itW8PHZ6oMLRU2Ak0SNG4f+
OKMVg/bCPtinO2CSWy2MoMXXimwt7OfkOtjiL+MrR9q38kMuj9JNuHXUPvH/pInd
o2cdI5X6bAvc+8/dOgaWuEwKZ2nk8nfscrwcc9fRgg9k/iJFEaQXEcsMpfpPZPKa
QezYrdnvIGbNkmLqgVYvcTEZni0LYhHZD4MBqDjshMsRfggEUx9L4aUVR+u7QE1h
N14k1juskwktw1qjn2p93cEzv/klSXcMjuyWChpUk83Qkxmo8FuypxBzxFEUDVf9
DdqwD2KQu5uzNST1f9I6RcBF6ibpijtHwyRJBptEVuJ64lwV6Oft2fobt77zVhse
bbUzA3U/D4t4XB1PNa/6ocd/AKg0tjZIwJJXfTq7xOcsqB+i4Nxh6ZdiCo17G5Sb
4ZrVtnDWt2jrqp5q2IjYDqROWElP86yaIH+2p2lZEHPm4wFdw7XsANgC+cZnc2Qv
69iX/G8EiofI+42POYT/kEJHuWmoRMRT80HsbXsTucw/G1c5O6x4sDCWYYoo1q9n
M4Y8PGZU4tgtlC2hR2raxulOpEti9JNvlRWhGaINc8pynHepJI1FCQsF2ohO1sVG
ZRtRn01dSpLRE8/8IoWFbBmHaEhEZLyOR6wVIkfODykbd+TMwilkEFjTnhdiOKUl
E6fDmRAzDfsveHQYonMxXrCNcVAPJrJMR0GFPZvE3YW8/H7mLDPV3rhTiQUOUvd4
VTvnRZgsrdLXKp5B/0Xt5vHm8sTyzY4aM5tnjdEJVR1o6nG7KsDCxI8GdrpMG0Rr
wV5sQEJS/xTZtg+YxQ3psIY8gTUrlYgYeSfh/rR/8kEDvWz/6TYqkFCWOZ+Ajo2v
8yYkOxp4wVABQzdF2/iVEn3Wd8jlbcNrcvqRsJWGgFh8whX8+s7yQIwic9anm1dB
HOQuU7CUDYwVOR2a7VXVeDw4008Rho28fwyGFryJAQgIhnl8BUfbrdV2vpgnqFAJ
DKmdWsKoQpDAdoaQcEMyUn2PEyTy4QbTRWDLPteA9+TSkWiarPTJtUknou+vSHnW
HIzphwUxfT1AhofeL0jVmwJYzk3C/ZMPU38ryJMPqUuAYcANgvoQKQkwVZpFTP9J
3DqdPl7GGNNPRJ01aCU6EngurRu2roSG9THvJISZDQEB/DqLmV7giRCAeDg8H3vk
YOQyBqm/ejPnXw3Hz2iWMLoJsA0YRNNAj5IQMie5Gy3sqtftE4Ax86WbS+CRbotH
SOtW4OmiF/rMT3ylKjFYnWLlMhvO9HJ+p3drtRhZpb1y232cS4Qkn9Ni+eEbzvL/
3FOr/CV/UHx/lw1GHVuXCrhV+XXVUb/7Ax1/M6vmcnh5PSiejZx90MHndpfYLSiP
vOmHSp7YDDfcS/mY6t5agC91AVwYZKMvzWuVbuOzvGhVyRJbNZG8njSGvpzsiabY
LJT18hsb7o7Z5aDlwE5pSwiWVzhHMSpAIq2ozBvZy2QvwWpmZSJMoY2pmZWOTkFw
iztLhwvexic7CgEu/+GHQRp2mjIVX6oa1025SrBq/m/3p3AkST3DmXgmu6OBVChU
ca91n7C+xIS7YTI1GvUxLlfI/8IIbdgsfkO9fnzvBQRSwQYg826aQ41HX1GVuBop
9vsCYNgS0zOsxRfCdODtolsR3EF8N3Fr9ms5To+JiYbcXdQWhEsaK1oDw7R1Fh9Q
WPy8v9H8L5Qx+6FKIs1VQ+w9RbdGEJ9UxdOuGlA9dJrOdAgaWKipOOsYw8LA5qxH
RMHjnV4uOhzL5Bitcu9sqLBYf4Dhp3fcRZu8QjJGm1sHP119SKYwk/rYNc1L04zM
Cu19OApY7yLqmEUDA/OOZX0OHh8tcuUic3Bk5IaHzOxkM3psj+rmxt4posDI4AS/
y4oN1LNtDzzbRjC4h5zxhWBpy1WkQNjq9+IxvabKsmQokca8KcFiHLWcfCsyURFm
xwuUYDLjio3cBmMUu4NDCxI3kaH3IAt+HH2CgNOriZ3z7HTr9Cly6AcYiOZAKc3P
S+6nMqkBWSfQhPQH0nPuSj50y040JGC71nxq/4wByxSmWlfnh25IeesJByDBQ8xo
HcSlYMCtQrrSta1Qg6uybygUvBcAUfUA+yUlWJcI8HOW3HkAvPqsq01KodRG8XIs
FO091S4hF6OKYDlG971LZDXXG4TWvDkJx8ErLk3PTqbKbk1eIjlwso8+S0uf4h/g
yT6PXBzuIEfiSjn4zdVYtbxRNYKh2afpTWw+QgC9bu+vQMi42Fx2QqeEnB6onuaf
yybaN0zNycX6wG+xFynvXN8SNev1neJTtzuXAEvPA3lFcDuBkWGia/sqt1C9vgG4
tS6GHukTT9wjy8wI5gD7Hm0SvM8kDcnvnEZMWI+IWm2WkS2dRcZBC7N3RBAMWXg2
IbKOZ9+w3hzuJR6Vv6qpVhoW2gAijgRl19m40IKcOjSWue4+RaGqDqddspqfeavV
W4eaaQ9r+0ksVjRO/dZX1MC/SJTsYno1ZENjuNAxmkKPT/W8l01AXGOGXnu4ekBM
tYv4yiD4G3+op65RAZXWmYHlMroGY+pSpx2Pn+lW3aq9mfMxA60ZqwRZaI6ydtN4
RVfjcDKL1O1oSo/gwKZxo+cQp8tusEOfVFAUw4kwVPLEb9ZHM5Qh/aa5vGRHbLmy
qg0rqbQJR0Or35pgwJpxQfr1U/6QH9grFmXNvYuiancbN4OnojLV9D4OJbmA9LC/
VsZ8qNYL0j48gz8RvHZ+PakRsJnIbXM1ZXs+/D9SfgwnapGzHT2XQ/S9NAMP28GA
RMi57JOByHbKQRIM4R5PIYSY4OLsxlGp++dOoEs504z0bkMRTQ5t+Bxw/X50CAtC
sW/9TUGZ1B1wNSOSilE04YVSB9xw8Vn/Ljd3tNPvj5zNqcDC3CFjjiBgghgj5EaN
OQYOQNDr1YoOGwTXJeEqxPl15hpxfS4tEBp80RF1fstxBmD0a++eSG4vvbcucmmC
gEK63XVFrLBLui5w5CNK4+wlShFHL01EEVOhrZCnuUbic/VOW8wkrmzYaqjuHPuR
zBmNauEAKxE1I7o4zoAUUdBsJzmVAet04rFsKVp4H99SicKW1atXbd5A4Bf+Tdb/
JiXt4gFsNTyv6/iZae13JTjiN92F+aJaav01mSW3Lj0CNRirFc7WJWyJ1mku7zco
dCfc+C9PZuotkDUx7qXsKr3dQxQDqH8Zp72UkgyJ8wujqtfhiA9vqk9DtAEkMKbd
C5xddPD5glI/S6nnTd+VZa4igZgMsLYm1hX4myNvV/3boPnJ2IPp2iJ1wheFHZAp
7/rzrjCncLbsUU3wdH9kKBW1HfxQGnfU/1ZQyafG2Ygk9qrO0SE28sna7xJnYdVe
3/ttZomldFs68RSmj7VeSy+79rEm5vPw22rRxiDPMz4vmmjNtLtoWUNQ9r1mc46X
IXKHk/XpH694LpTbKqwAWjogSLrBZM7oTNGdJf9lo59+XzKyUWO09Kwtp8nHEWV7
rE5lB1QjQVNnU/bvzOiyVTAMPq63+se23ESxdj963gzDimZN9y0xEyOGFxY3YryH
3Ux0x7V4dieocoFFaYXKunKV950WhopUzCh7r5bccOtPydSkjJ/zYsdOhBlzLrPX
Z7f/QBvZBT4HsER8t31s3jAlKqZdlADEraL8g7MLhIjlqS9LV1LIFXuvxuHvYfhe
BK0kbyWn4mEoRlPuq5YakgKS8/diduJUX7yMl4x8g5IqnDrK7IdGVRIn23V8lWua
SbB2XBoUbg8p1O2q9wnxq33cMnvVHpxZpJ5LbiT012zL3B+YPauyuACj1ceHZtKT
iszvyvK6GrlUynVCL6HJQvjNOO6l4tTCLPlW9ilJk0wCLUXHYn5Y+1f+5k8b2sPe
yyCs9cHZZIv4Wk8ch5UwvFnoK52bMKGK8F+ggJcjSZDuzyzf38s4Z1huhB29Xc8/
yB2tuHaH0ZdjdzjN9Tid1HBNGEhbT2Wm1ONrNthULJ28STLCJlyssjigqTPNNmvS
aWAZDMfM2k/sKYnUwfwSeoL2EiMajQe0fdwOG022B5wjtBYUBSRjuVBzlpbwP5YG
+u1hcYrN5WgKvXU9XhqSmLkonP7/1vhekiMEOgHH1/HyufROPBSno7J2ZeuyVFRU
8L0Eh6JhziPUdhLt4NDbogNrksUawa6jBzuItw+gSiZRoAWxHfBZbfthi29pZ6ou
L8tQkr1bn7hvA3HRKvchyMx+W3ELocXXKjKWlywaPVChtewtAi2/6HFGi0xyruD4
4MSj1zFaJwIeIe38WDqoDQeP/MyYkoFp22truocKYUukG3zVK5DLRXf+zZqlkNds
8KqDlcRVfjDyymSng5AfwIgPxb65H2ekBPB96Nt5m6oe9urHcS9pPZ8e6wobNJ5+
o/0+Jy/VENIzCZepWyKLVFPyp4TesqcfKj8M+9E8cPioJemnVgPMqxNdl9GOeogq
G98lFd/zbG+9IdGhQKGGHplC2oiJDEmHybySv7F37qvE6QnE1kMn3iMv3AXbseod
KIKl2Ox70xHA/aiHP7bM6nXI8DmJv6mbdfaWu1wV5ENz121AgLTnn4p84u0WqBqK
w8nqN0XN6FqQf9R5G+KY/5wxsaIChOVgQUJb74GeTMBu0OKd2JzY0b6dwjAAaES1
OAXWlXqaE8lMtHTtpkHgZUCgJxQTyZiMpXvUVLXL73Z+DNVaX4i8Kf2FExaFR6U9
CbuYYkzjLDkdwtmge2RHlTa1Z25kvGkSKwJL1IgwV8N+knV7ybv1slkCxU+38rMc
BThCqstLIRD+mGhzSwCULMHna4tdlagBguiMmDrYkzOvTEbnGtgU1M7AFjTNrC+d
le0EZGYctFX2YiyN6nG+177zcul8ILSIAA6wIxyD3W/sYhPJewPa1boLg2l5/P/g
zFg9s3tVpslXaTkaJV7R2kODEL3CQpcpyih3YCNowUKPTUNoXYt9k7WFqrbevhal
6wCyv4hk8lsaKcLfeV0NkoWm8xtQW1dVpbE4PUCEfmTJlJML8xNsEcHWa9U3viFu
wfVL2DHqWkO9RZ1v/d3GCC5k/kSrvkSExbgMWz4xbnVxRWP4+miIlPvCeSvZmFRn
gXIcd74H0AHrc9gP2dCHv2AGnjjqy4xH1fim8Wd1kpXEriT0GSHo/TV3yy1TNzlz
l+uJ3wcqPle8YoR1tf2mj1uVPI+hgI4tVdu3IYGKnQO14KgqDAjPkytkXegEecKc
TeAG2q/LJwS6DHHnNgnhwkSDu0oNAq53uTCAVC6qbEvw4jypIecfOKJZM/s/RUTy
DfJaU8b29gkyVC2FhPgzpWvvH9PPQMyeA4mCgAK22N3sCot1PgYvF2ksVgGRq8eL
oQ2ruOTzjKgagv6FTI7moyxvenzbQlqlDfgjgKbimQQXmXcmrEc96d6KKhmswZb6
vC8xxo4/eenxMUAjzLdJMCzU2BZPDlp9qfDlw6OZblZCExOAtDLW65TwiruHGEPX
Rz7PJSrZ0oEXUkkWNCSPMIoTqloq3XMA99Wq9ZjBnTQFSBrFpxaTFhOcjRGjRqT6
oIPy09caA835uQBib8TnRk9aeTruOqOu1dMJ8s9jsVUCVqMZuxLPWaZGtLIDQKa1
1CcuPvG8Wymp1fvYpd+QEn3xILKyZURHTEA87vWH4RLNtsJ4LuWoQnWgLW5sX9AD
Uhmfo9qcAB86jChAkX+G2eDaSSaAbEwCoz2DT/7oPxHZt1sAYPDodoYuPAXNKhFv
3sr/IetSwPGgWu0+/EtQF2cqwW48IxLHU1Qe31CLKzObNrwEuog/u/h3roMKSQKV
cKquz93d0zj2UaXWUmgJdv20FlfmCiZeul3zGSp1hQwZ6ZF6mLi/nKJMVP2nLRHA
jUHqVarIvxIrK3JDWIJBlOUvjyCBu3hBjqE4T52HelW4zI+/d69j8C0um8NHogWt
xq9ch+LWfL7AWdIcA7gBw8/BSjKTbeAzuspFzY6eObgDPca7yu9RfYAyV3tpYoGl
6NBfWxvqcALhwOUH6eW7S9zKED5IAYSiFLJY9c8JwFTPWI9I5/QVScxeUjE6Rsce
8mOsALJhl1ogbQuMuQWGA0+/k0tNXelxdvHqCc6iw1fCDpX60tZV48tue7B3bgSJ
aFr0eduNAsoHu58nbiSW8jm+EJ8Vkbd4b9ILYuxqYG3Pk7GC4jQTIeZSRI/ubdGe
myzGfbR6dOnJvPSPQf8CFS53adswtKwap8wRnrKzkljlxhzANwReoBRtyHsXfobm
prjU4S+E+kfDDNSKiMtYshnXR1imPJ/OkL3Q6mwgmwPbtFrZYaX9YHNVThVOdSz7
djuGJ2gO1Hhz3HtJvM9FCZ25GUbies0+NwWyhrhKxizpCeXAbsZ3yW7J+6H6P0Ki
YjLb0DjoMY97ANsvXW7cNJoQFcRIyamTS253D/CsKXuaLyesIfQarmkYEyoOhM93
PB8gzUzXp5M+mX6FujjHOBgHvN/Cztd/rS0pWgVc0k6JXMUricyutHuv6apOAzDH
e5Px8Jat5RYnTdAh9kulHmQpXghNuz7GUIvicN6ED0x0FB4ZsXQz2LU7RSieSAt9
+5y5sUe73Fx6nhK4B02m9mj1XeFvIt9FJctxEYYGEX7HdpWT3ZecNZ0zcV4mL6Lw
SfGxrHXVz/BKeRERKF0Kp6BW42g22Z3nriuydI7+48N6DK/bGFDcZqZEEVLUPRPv
4tpk3PT6LU7eiktXFKaw5X6F3xpKE6WKM8nN+PEHmUPB6Jg5BdZ/EXQ0LzjyXYT+
lX0rCnzExCbuLBvkLl0in6DpX/GwhSFzcY1UFAOGmw+1WBEVkNYzeXVZI0yMViel
fgxvWoyFL8fyMWZYLykzWY7WenwKqItSEToSBC+96WoKpsO/XfmlXRqj7SziiIKm
RV59q6yoEXkyMBFh7RgaZri6c/unmC8IP4rHB/hj/R6JtaGvCMrx6HO95UYJ2Cf6
aK29C3uj475pUcFibT4CGboVtcBMSeuCG3dsqPw+hXwZV9v5RZbsV4pGGFwW8WUx
Iml5kG/5dSPqGN7E15UpMGB8Y4JlMWSdMLmTN/Ini83V9h9bbiL/U7TijZdlHhzt
utHeJW38zV1u4Hr8zQV2LhnDtHd6H5J6rC87IKe1lJNNPFMx9mgCZAwxewc9/Rv7
QOBWo2YWlhPFaGlCpeFvRmI7JxMr/XCeDAdvUrLGo9DuSYqMZy0trmlRIy4sHoyl
xHU8+ZxHpPclqizPFUsqjomM576cuWUIPAo32NF05IhYnIyIKtITwaf73CLzX01Z
oRwtBkVwwIcNZWRGT0BQPdMIJAgyxqRRGmFcsaA1FRZzEAc7aJ/swO+clMBLNx/w
XCgfgtxEdP4TO2n86hFIaPoJpRAodiXRzZvUmWb5u8XVg5XTM4qtifGF0bZ1YOVi
rpuM5HYPhBiGv+Ikdm49A7dmgpRkCnxIoCb5UYc6IVr/XH2PLqeTn4vvSO2te1YN
cN1jVIttvCfoQfQRkC3qepjjbUq5lJNvexY4UV9VsaX3KjSvqLzXMN1R1of44lGj
A002DoCqPG6xXuvEVNUfvQdz1WPrqluJDVXrXWrZzLj+0HcCneoRnpUxdvQpOMbj
DNxuxTYy55/c+m9ZZHPjXFk+1gVCMRMUxB+jufSFlezvr5e79qCdm8Wx0bw14+Vx
KGm/xTBCVXGjxw+Z8Ha+OI5FELulX8FqtrBRR6EQFI62XO8vQvWGpsTeSTNBVsxl
ZpjD/fhcU5IFJAh0X1eO/BOKLJmWqwPa+9QgcHGsZ3Xh9ip/2jE7ZtM4Hwg3mj+L
0Uh+8hsNsa77UT0Ay7Zb+Q5dX1rFJ332J/w7brEO+w0NgSsmaEuzh4z0Z0hlvOfo
BuqJmpKE0wkCWv9rOu0DfhmCBhHgSmgDSwE4WhJWBhCC6y527l2R2ShdX6NFhBCf
nMw/8YDCQS3eEqjrQp3VU1ER1zq9O6PRqZg0niOPs4kDIHq72KNGX+drr8b0lwRW
8JTxoCqcqxWS0P8Qp5P+nYGR/rO67D0CaFaQwu0lXVL3uucRferWqIJ8C0Avttr1
cR+vzMWDcN3/8KClamEvu7YYjTDhSpetMrIxjmmNXAnkoyJLydi/wHoJ/Xfgp3/Y
PYdOSE+zCAjjWQo5jOW2tXGapdLIsyCyeAaTQVEq9t8G7OYPzyegLQPKw4kCicx0
hX/r+LL/ZdtiOvwjUoAPzFCYWoaege73ApYRmoKTWUcCaUXJPEdv1KYXvxFHo+XR
j8DOvMmHESoCM48Ut6P1jVjABXQ0C5U2SqsWnZ+/pJkP1ZNyRDeYZGuydZ6d9sqi
AqMUt28bn8cKs4Wr8yNfsF/EDSrEaZn7yDhjeMh8qe7K20G2KtvSiYTWgyFwTVty
3LRAbaWfR7gHti4qrN1+O30qWe4cgLKmjswv08/4X5OQnQKxtazQCjjuo3la+gvt
nosqfP1U/2RPfCx3FN32WxlrrlOL8x+sjaCujsVuG9/18ZHEPO4yOPNUfWzUYoTZ
I3VmJqNjilVZ7FJGWGrydYFTSJAKeoypR21Q+cvac4BM253+rkM21nEJxIQpff4K
cIzzvvUSSP/fO1toXnBlE5A1/ndUwm0BkVvrGRI2sUY+/ySr3CgiayyWvXbrNbbu
SPTIoXm5cet5sxDT0Slmu7gVkypeA2Xq+G+P7yPv1dantkFH7X3bq4/X+SM7AHlj
IgLMcXK+C1dBoObZcIEyDDfS/h7LVdf8sHa9dnKpKp9qyqKYthso/9vztPeUBLsd
AU5XJRM/QUlp4zVx1Kc27B+8GITnM3JQyBUDEJ7kF543MGuKKTBvx+cLYVk8a4uu
19cy2MXhW/gDj4qiEtUYpAopap8dj7zazXKHNhGz64Uca8Cq5JyoTfu2Nivr7oIW
nmD1/CCrr2k99ZbZvxKgO5Xr1rMg1OY1fVLTXiYTVwQ2Jn19UoWH92W3tk3Wp0JE
Q+ZKeuniEslIx7S1OiCsYmxoYtW/6d/2LS7t2DzLepyEjiWV/RZNGGUg7KPaS2dk
2BiB6Oh9CnL7VMCn4sS+UF7M2uAMflbJVT5rqZOpxDTtXPyyscXxUdFS3VwfFrwG
ibRcRhoCy4qu3n/ZwuxHiGnqdeNaIwKSu2Gr2q6dGs/RGPKW4pDtRCmZpj6VLsbc
9sVMoh5ZCZa4pEPSSH0o9XIiLjTCNiIyigEJjGQPGZUeNW/Vf0iR9p9GObAbEdnL
fFG6t74NuHbEIWipBsAihIQC2u2Kx8bUhOU8N1qmC3CVU2mE9WQMdCNwJQa0TSXn
KpKmZeSY3khQpwlsfQa0fD/xfECmLufZj8VWVXNcpZ8EE3+ICtY3TUwuJFcwAlI4
+SRjM0yWMdTLQQDnB5CfgURFOgF83Va19RbZSz571JkDyIlygYdde+LL2IQxTDl5
2XgnAs6eKc1LBgSjpUYjE+016SK3E2lkDoNAJGYA4e4SG6+ZowIQYxXubuPfSYpS
iEzMRlbwTqIuYZKjMiObRMxjtHNxkwiiNc3zZkHUcriaNchxoryPRxCd1iGGlXZq
YN/feQLwQefznOiEd5NUf7zB/ecTV7dPBneOASCkGPCUWnfJRg9lLT6r879mxfXF
XgmbOPQ9eDCeJBLFsNBelI8BBrTPEvtFzRbNsSYiwWwYkJ8a4ZvdpCc4RtSQbbmv
ONe21j2AYL+FP/j33N1H/y+74o/9Y60sk60KLVGY4IszD5UizGTJitYAE+5LG0XK
yY+fuYHH3XPO2zVTewvtPk3xilQw1vsUbP04noE5+g8qqKNPed4q6AU8ZssxWwyB
KCYnyFk5o9bHOwU2CF+n4uyp6AvLKZx0hIu+9ODtzAJRaQyn5wasH/m4ChQNN3Ws
c7ATlPmbvqerOhPA0nTWAdD1v1DgSzw6u9r4MuIlMLEr0UqV8gwTpYR/K7PNiEk4
lNnGu8v9i+oyw78A8nbee2V1VI4XjM0oOIRSN6oDvQEj5bAPJ995B1isN5xnjrRE
Qb8kvvVUdSg76e407WKttUPcEpV0dn/ruFScKF2ApEtJ3GptmkcU92h+Shypv1QS
75xk5i9tqOf3lXFo1FHKLGvjaGqDnu2Kic3UJbNUlnmH1ss3m5mZdcQtiA+y80bF
w6ZYXSGC9/TMr0qrLX2aOoRTur4FWDh0n29j1xfFPBcn5YUkoMJtWArR2P7l+Zfk
eVA6Ut50xczltVNVe4xouSG/EaKoBUnMH7nbrNjZ0DYDYtmCkNXK6iPp8DAv6jOg
UqlJAF2XHtRjdt5Xekurp94tM6iBPo9qeLasDgv7ae5+y3Cl4M9xn49FmOGW6ENr
2p2kEJE0KgitGSdwHLPqM2bb3l/TI9cTgVUHyPwSe/nRR6A5ujXQKMw9YP0PFFl8
yye8CA1pu+QnWrc0i3laG7Q3rfnsu+y5Jv6PQxV8KzPniCQxbdTd0qzYokw2CV3h
A0Mn+tB1ePy2mg9O7+FJdJ8XOggUUsoxdPfiXfGcnnZU4rgRTY6KVS5Nb3rnlB37
jaPVARTL70wBXHcM5YrpRMcrrw35aApXKKdD21VtqeiBz02HdPDlPEW+a9a79Bwu
0d4IVQbYUsPkLey77L5m713cWOnxGoKj3/UCXs7TGwvbrTH/EuSkfX/dQqkyOIV4
Nv6hGIVLJuMIPuFevPdUt4+dYHQPIBUdlNxjGuRfVapF8SrHgjv7HtlU4bPRsE4S
AxDdDW6yI3OFp70pzHwix4f2XY/+6erbu0m6zdtbOZQsXyZV3jDnYEqVDDfB9HUX
+TE221DPC2joSZb/GuP3OCKGS6gxu4lauTo9mMboCJ/ohL6RMFgPfuRXXl/Okugw
+nfZCkm6lUoP54lGw/9WRm4Xb4AdMdJvpeaPSXZ3TXMhiTmFpDm1N80tAwl0lnYL
oexEaTxkvRsORicZ+NkzpfEpomDyWzS+vsqlGvReM9w9L4OdzQ3zryGURJ+2GJSx
unbk7LZqdO+Os9tmdqbsp3DmJvPebXacu2+rGPwa13XxRtl2sMKspZyOIGH037ht
Eqk4wyag5oDkoMM/gjeFftfueqqQxndFIh1300vIt5d/K9lKEvE+84RcGOuwOT3q
uRcm8Y4MIw7vrpIXRNFaalCrzoZXzRZsrMafoTQxdHpiBBWVyo3pCfqQz34kO6SI
DPi7eaOkJxU2ohklM8edqZeCmCzrB2ezQAEdHrSWtzpyVPc5tEGW5s5au5Tk9uZF
Im4mfs3MYzojejgqXy+Y5ye+F0q0ni1EScBNMZ87fLPA1AjpOEL0OVGCOSx1BDVQ
mFZ8/kRpy020LRQemGonmHDlhsWPGLbvYILS1lNox9uFGKZ4P+TTtLrwveVYNjAz
ZAF5mQ7wHBurgTLMwU93xzfZrj5P6cMBxcyX9q966197mA2cRIWWcpfOTWekivPu
sdNKllF+hxXkU7hLetGv5B4wasK+j+1/e7ZAR3KXncx2xA31Q04pngTzKAqoeLZS
U4gjEHJcsGM3Y/EKubwwqtjRToXksbAcISvKK4Y2EHKr1lGYspJO5cOMem0Re19U
XQiBdTXKOn7g+4TjS3tdFNjth0OLx25lKcuH41UvAw1aPzVyP+8CkxDIcb+Pk2vP
6D4JZwRpemQoMH3Z0OoJXut4dlUjUy8zq3fj4jvhXUwXz3PI9DnEjmZlGIsk+uvx
MFU3H/TvTvyiGrLxNwqYhFd1k3pgNLyVj8XDaPN6NtiB1tDFTUr2X2TZjO7z+Rzw
+UqobwPbRx+pWCmEswK2e5opWacUvwNaaDvOs3muauKtdW0du4Y8ArhPA0uwQswo
ZculeQa780RJxcMP6Ed4krN7V7KWhbZE4SLyP5QoYW7slVqKyK/yD6QXBizb6erq
JVtm8mwtzmXCOHbqijQC9Q/QhLe997q09iCbysnc7Rs3pMrP689KFlKhgg7youZG
JenVgK8jK6pOLTGZAqYPy5TgbgNZjwf3eYzkdLSWP6BH6vj4VQFnqNrh9RSrBKud
PVaNC8JN24xZ7wZk6ckgcqwZ15LUtgIZ6zMEIVGdf3yIZPuWr9lKZXasT0JjuNuL
/TIzJDYJtvy0vA/s5++0tgqVnl9jWkPPIMPjpRUE+pPQ6S/An5qpskqebbb33EMf
7o7hkwh7a6vQ1iK+O6y3HLa6kU6ZmaQtOWu+8GQrWOQzSbiR81ic5hC5LEkvP4Ij
i30IzgQFADhehI+VErCkKf+7adVq5G4GJH4b1O5ZQXUw7t11fVycE4+FUABki48R
Mc6a2aco3/24pxK5Nbsqgw1bypt1soCR+3z/Jp6eWxTLmEqQQtcCi05Zh9N8amlR
cX+poYY+vRW56lp805UBvXbPT0RBMuUUAQpu19vekghD0bXO2woPyr5J6EMUQTde
4upUHmMYo1wP44+6aX3pIP9Ykqdi5zopRJtDxTbbYTxQp48Skz4N53VHCoMTGr7Y
RVfGjGDWvUBNmzdxEKcZf6ipL7YSS2uGeIhwzICvqsQWYKHdS75GtJ/itwpc2Xvz
I3TlfPOtLoJhPekOFSVsGHNVaFbXIWT3Ut/40kHrkSuEf7oEJ8LfximTPLuLld3k
XCokB8tMCmhY8YFlCk5z1QYC7K977XF8DQYkVEJkUvIIxaWY07i1MgNBFWKPmMc8
UBEpZ0mI5IXyaVmlPWS829s72dcSekLkAcjMVuLHCBjWAQI+vUE+vCen8Dtgb+k9
E+74NJRqn7SGkMFbOnq71P9BfcDOpPDSdmoIB1NtNL4OGqyka/nv83wzA++EMeHt
MUGCFWWGDBJGrp1eqHkFTITo9JojkozCsMPj8xbC/ZJkmzJ1yvYQHmoMWBmQNe0H
`pragma protect end_protected
