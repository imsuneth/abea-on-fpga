// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:06:47 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kG/yBgigY/LSaYDue/n7X9O7UvsJoTjpu+81UWwoYBSg5c3tQ4UPTNuGcCVSKHeq
nhR8sBGLsjN2Zc/4R57j1+d5sNPWA6kFnSwJ8O+j3SNEzfL76TcF18o/ddaSMHpZ
tw/g1dSgeZIfcxTTnRnX17rMTE5JQ65AXDaKGvPOr40=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8384)
j8li1KRTCT46J5wW1LDsq3Mo6B4+qphKvz71rhg4+JiLpc1iF1ccv0FGzGn3LvsP
E/6IN0aasjvaxx6iVfoNdU21+h0c/H6Wk7a43OCqC+UpDOsG5Ay+9sQBLIkLJRcL
xmfpKagmL17scCGWtGoSuv4+AqPHCEmWct33NxGpCT7ik0EaQ42w1M2GkK6Y98eF
OZ61JT3NyJHiWRkiMddN+12RXJk5Mzzr51gA5FjT34K8iU3B/qcceLfVOXplhe1/
MeJsT37TLi6zn4lS8aCp4gxFqPr6YLhBWNV8ZBXdae3WglvIyqaferSNCNWQEpiG
vT4JtB/iRFgmYxR4BeTMn3eNN34VzIFkYrTWl8u322RSdb0MXJvCdXNHlc5xyYkW
T08PB7YU1XZgWnlkyNOm+ogeWiNKS6pPdWy8ruBADBBjiYCXkVQ/EJ+RTohyWXqg
FUHTGIPfZ0GY9LWZQlG1nqrUKKm46rjg2uBLWiN2w6rf8c+dFbLbaxHrk1ZW2bdf
exvByH1Cm/6JrRLn96u3LArIZP/WmPmLv5B/2lzyCFBd+RKIihAzcLbPLldCxMdN
heULQDn5xbFGoax4vGhpshc31AO+mFWjT1s1GyMIhlhqferJzOUfTd9Jeak4Bvvt
XN/CfZvUHvFjLBcILBvPvv7bNUk5D3qdljyCsmCWk50jX4kdI5XVFRSpczL4yHe9
hgTo15HbvltktEUGbZ+kj0mWyZAxdPygdQhFbUZdz/H4MmKRY7aXIFUudZEoqCJ2
iX9sxNEFnrUZ3HabkeiI2QKwU21iQ8jOcsSDKyJERrr2dsFu7wbvLQdO6rzSOX/i
Q53RHRrRb4K9qoqGkfdFIVlXIUwtO6q9q36yEi/vspY5mH9c5sXSajts1hJWjDa9
0DyqzZ+TdJAxJEOCiytDrn+OVKBQPPX+ia7j4ASghDnN9gjXOoBAEAp07FACWa0I
KoPgOlg7KflI6nWs3S4cicuHOKyLd8DDcIPUhLZ4AGuves/lLdOhWK5s3PSecDio
x9lhDC+eQweUH6hakNGaw477TbwUM9g6yYW86s5NVmMucwyXZXzaHp+v4cfXdkiy
G5jucFQ0fX9y2P4PU30iQ1SZcufXePUAIxCJjoNdnp63aJEHBLZypoOIJL5VFhiq
E573uTGrVSTAHv58+IYflDvYs7ERk4WizYbAAyshlnrurC2QcEtzLMrd2T5X/4Ss
660QIQPiD66kzj9+8mMDKDxfHyIi9/169m7K5P+XphHmdU/X45oeWVUCX50RC5Ry
V8dborbelVi663BVO7jjbnieYvk3EwZnee6PVQ8scNkO3bK+6LKmt2zPZOZp3htl
yepBuEc8UzRDrUbJxnfQqq0DFL9V8fe3H4BxgEwF1TMY1uEmdsSkvftGv20RieFJ
5ZiEAuEVebXi0Iguq+q5cGvBQoebjJya6nVcU3abF/SyWj/xy5hwCoQRUJ9MTdtH
A/t9Bjpm+WK9C2hCfbQAiMsmJzqwnf/cir/8sQEfdx0KFIa8ekd/3gePQYwhAoIp
+5LQ58iHJW00CL/1NdPMU7jMr+6DTQOYrCv/BI1a7d8wkNcP24wBcTiFUSM0cTxy
cyQkrd1EZ237fK+TaQtUWiSbiYktTRLeZ4STwIaYeyirMrlQiKdYFkmj9X2aH0V8
pfOnPr9kyQmCpJcVUQoh1L/iP7Pvo3CQr1pNnlpdb4NRjk7idTt1Cctu/C9T478v
26vfzfCNBLbD+KR3otxUZ01WGUs6Tsjoe88kx5a44APB2pAIktyb8b23mQCTlRD9
Pref4ZS3oNIG1/ilX80A6fWC9ChbUaMjKw1oylAxuuTw1iI//5heIStMSnqkj94b
qdGl+ksBiCSs9Z+p/+6+swB+KQvFTcVwSb88ovYrtZzWhao+gqCLxEfaZhf2Yum/
92QLKOvhTupHWwb0VsSwsjYjEuNPguTBjpX1iMKlLtNtwqn+awA6ErYgXq1Iak5Q
RxDCi5O/558V2Rfh/+mRiaNEsicwdgZXRUOh3ZNCbx5LKfszTPzEGvhtK7TYHSs6
D+6dFUMNt2liKCpD8gl9vdkmP/QTN1i5t1rn1yrLvep/1cm1dg9lADd5GPSBUmhI
XfN9+QCHc949U21pQLjfYK4+cwyuyXDiIHzxnz4mTLGMBcMqRlZCdwVJo4TFFRkJ
L4EEMgCWqbcNVbfOtwjny8RiBFtdWq5Zl2VzZlXhieFA3yjPwGMOLucoq/9LWxWv
8p221hzG7m5B4LmzbJViiy2ISQobbZ2orpGDCvPQjejSqL2YV/J5mtkDb3ufqyjF
f9+J2NL9emVFC5or/9uh/vlukiw9+qKVFp58+fruswexoeBMVYIypsJJYQ7TdEy0
2bYiWqngy+0elvNL2rovgXadvTZMR1Pp0rQeDrrNLGBaPVxSisK2wKkSzRIzZEz5
SYlHxm0lNYnDYIltCycRNu1hB7QsAv726ZhH0FcsJVNYwKgjKe/efirpuHfs4ZrO
0FLVMYuXmRZgk28h5D9ngt53DTBePlitL0hqs5JRxOFW5I24G5ZKHO2lcjQjPn84
63HyGU5K4KRjP/5b7Ln91jRQPOulOmxuu23m6vdeOj/l+M9J3DtVbWdSX5LCJaTa
M9hLVt7lCvatKKcyr0IbWBWqusAWaC/0Q9d4Q+8xgS+H0yvdgg9ICB576XuVho8U
V5l/pbVheGZgDplGAA+6+kBa49qmrF3wvA4S+rPUVEQFAbRNp/uVp2PNTWW/w/tJ
DHBflvaOwDD4SJ8KFR0LMD8dzMKuJgkIRmgDuTe5wtVdhpgnYZIsyEMlX2lGcnD0
SlRPZ8wE35RW6M8HjJO9uThsDYI9tkNsx80wWi6EiMVBtZpUG49nxx0xOLHaUZiz
+RUhj17wjDrfAUJUiAYSu6u6ut+h68pY7kSwv4vQT/kg/n25MMK0iefU5tAUk0m2
cXZ1IdZNd9aNNX0aYSB9vENDGYn0rnkiFQPjq2JXCt1cO9WAU2o4N4yjYFPadlCZ
FQhKDFtEjPKryOvPO3EcbUt6epbXfjSXlx4C+6kak3mQuEByMyir/a5UWiED6+ah
PSf1eoS3LzG1yFtLzqtcl40GbLfPHEmb3Kt3T6BhqLL52+UYjLlwFr4XU8+vg+KS
MCQtCav8RYGxQiqmXp+yZtVl0w1sBqxo1jRZaWvFWXksBmGZYCkRVC64szF7AhKD
a6ZL5Hfbgf/EbPQ7w+M/MU8rw6F52c34X/Tyz+Put0Q78Qit5exWP5CcRKnm+Gwl
oesmbfCnIweCYxfpXwoPliVncLBoAJoFVDEv0EH1u2X2/93//H62GSIVrNTNr0Y/
aznIwR+Q9vmSSjkjjsevxu5iywZhRM1IwmSn8t3CuPaTua4uY/0/fciaVwjifaFM
gBHjxkzV/tp/6wttBPqYphxrLho1VFYGMADYg6r+VFFLsm0vgxWD78HDDOaP6ggJ
Wq/k3ry6CNBIS+Bg8QRJqoPrRVjOWIy1kaTjTKgEPNPR3U/ln/na2fCnjSNwOW7N
K1k/kAUUs/o0vRuMRpZq4kaJYyEEZftrAc9qsSVAUuhF3GgGBE0O4zk8YdIQDSd6
M6rhGSsstcIIOCPqu41MdQyxuDpoENZLqU93nmwSdd91f580yxbuboaN/msAxl2W
16cA8VF5Yz9x76D+sRoAsesQrqXM5ix6ZkGfETZYu19eHC0GzAg+WmWX9RQ0JBgM
BdZvNqwsexaQUYKT+pUfq5BfmKUSbX2+3geDoazgRPphVuLu5nGl6JXmA6T63aH/
0t5fFb1QpRUolC8x+AlPTqXmjnOWpYzBaml6XLTI9Rxcxl1+t91OowDyqwcwz5c9
cQ6v0cLqckk6tZRFz4A66GOQdEDNBZgh4PatbKnTmtvXd1zJyadB+aLQlBipQ+36
LnJgOLq2fXYJxjnmE3UdHu+oc4Ma18e8YT2LtNwzfP1+h3Kux/ujzEsWTkfAvHvW
SSwP0pfVSoCo3jFwMv3cIDfHrZ0iDBFUQwvRSzsMCrDvSRN9HCW4iADY7NHHAXjv
QIpGcKNcylnU6GWq7RJrZEoUOdHDB4Ue0U7PH8BItp0TK8TTxl7Ou7y7nYeVZPJB
Be0xP1bA/bj8kNeyz4zSKzTLI+pSMvrsdbCPRBnlrhQ1KVgMN7Tk4O8M7Jwt3CNt
F2xx/rd8ZmGvVmXu2tlbsOkPAeEDsmgzUB6uIpwxNhFUOKKs9Bixw9LXKXrovMzB
rmRKv8/CQegmqR2TFefX9DbwfSrwEps1hm+Ga4RhrtvdxkUSwzlIkKrap4Ihdbyp
DU9AZ0vg6mn3RX5F1/wHayqnS/9cjeIdZoVtQIWX6sbhvpoNbo1jeRXt3EdDrlFC
DzmlQdmkBxzIaxO3dcHVpx7p0s/stDw+eo6hoFmBwlqrxlXbEFLVQ05EOwkNkBiJ
xPz5w3h4V2iT2U5zMRdu9hEKeGRhCzLJXrbCiErFzylCz8M3D+fcyZKYFCiGKgkK
7CjIC28BTd+uzevY/qeTX07W7H0oRvz6BMaN7YZQfDGvFwLLlv49OnbGdpx4pH7I
hI+U4+2E8JseX2w5wQ9puAB6wVwlF0xeNc1ScjnNueO9Xa+okKQQp3UBGyDmxaH6
enVRm4PJPgfEtonF79kZtbYYfdaB4JfhViJME/M8HFCZzcW0t1LV+t0EJ/c0PKfQ
X8DAITBbZMBq3O4wTfshfHXTsA2kBnhTkQQmOcKba+AWEi+PcD9Y0vUIiar/Vgik
l5CELsLJSGHRmbe6vv+TnQQp3kCaZL8X73UtQKE9JNaVwHAcoGHzD/FT6b4XhMPK
0QJAGVDaMqoQ5aX7wvs7gyzoYigvitsTnCbpC24CKFq896T2HUKrRYK23IIs4DYT
+iELjDX74FNW3IV92ib260l2u9kZO0VmJNEgDVainHbprT2a/bEzaLKeHiIo6bDr
1pNZPclY+3GRdXKwNdhyJQbJ8OS71Y1Ji1THma8dn+ieJWUOiTLX/apZleoJo5fw
dZj84i4JIdkVpHDm4yNKvPx7ToQyzZLfn8idoRnhMkXqbyo6zB6YmpkqjhJIbw1R
P3QBT2rgoSbimjJJ2xasE+5Y0RSm+ttlRvBC7FpdnPSoPzJQjcS31el3zi/0IXky
j4fj6YbaKRWVpnfd/UKmTnjEh6cEQurTFGikn12Bw7HtU+XsVTWZQNnT4Ss/VOLI
czZjjOk0ejiK/yqpsNpFMqXvRvAW3nKbZA5wFHJ883+nn51dgAAsPg0p9SWqcnU5
tUY3ao+Ui/ma2qVdvuDzg3IYkx5w5O6l3GjFgizjkbVjT+lOT/mRnq3clgLimL6M
2S6Nn9/9AgXu1m97e7iKn12p89cA7dhfyXWxZrfrACl5LOFsIlmlRG6oOamMRgDh
97RxvHl0y8cI8R9bj4FXfgiG1i5vzm9kSlJrD6ZDJqgaRe6XyMVOsHqtanqPM0mn
0fO3nvRWZpewYHsrnlCNPyShGlO8fd2E02pSZSIjQ8dSCP+xUL6Ann9rPs8av3fc
so1zbHLWiRwkZgiXDY756ebcZfpCp6d7Hski6wT44ZQD18UCf0wTGsncT0GgEmIU
maCMvA5YwxIgxox8QyUJ1Keui+qzl7ac2cynXNdGYxg2au01psQWVupMMR2jnFhR
9rLyg1QsIudo215tUap6m/av6I29jEeb+Br/NfGR4hbfGgx97N51+BNLfnEcjYAs
mb+SyyLeZtx0xrVJ46g3v9BNR+tg0wnAEXFrmX16XYXdR9ozHqxsfsdrugpmqB3Z
fyMTesJ38hLJWPDHsQVebITqn1BNNL2htFCcOfMyOLT6JVqFb3eFfxDfDgyP4e1e
1uGU7EYO3wMg7EJZa7QgJlGcZ0sygjxaqOjhsnRHXWTZ8M3JfepYKUtm7GHxp10x
vJMyQfi8AAE3awgbobgmA8emHkjmLHyDDv2KrlFvJk+V8rf7tMpIJ8aFrCZ79Zmc
pjbhVzsv2fHtPmCFyZq+Cmgx7iw/+gskWOjZ61PaWi//o2XyhQ+my8QIWvY4TfVL
vIpEu57/rbbG4aQZ/AD4H3tmjmh2KCc2zZ5lez8Ou5g9rTCXMRbA8sNisEgX/N29
Ot1PlVBreYULSMQZtS+/OkwomC5nBS7DDKoOFadNCID1Q5X4asCv/eU3Md8pSY0b
vwriFztXVZugSSmEkZT3IfdmhsaSxJMjkhypZ2r2MFQOb9hTM6Wy6JxrL3Cs92J+
5Q/l2XrF9iPY1n/5qKHRDwG+iBlc8gkWgREfWnP97hks2wobHScDKo4/qtZN8h6x
RS8YnAHJt4/8ucI+v3zWCITbbvvBCCNETL7Qu3n6Jf5wlSx9sQ0pDet47LuFpRnE
Wp1ntsOWEn8s3a34yW+qAKH0K0X1VgL82TUUfSGsTNgOBS8nOeYzAFNEZYQJO5dP
8eMEH1s7DgAkvOvtHtrSdbZhTvgcPpQLbIqYxvTqm9hOKzGG26z+zUOZegvDUuYz
CU18P61xgfM9VGzNLribVDq2xm2pAIcR9MjhFjwTg7taiaE6LpKzz3GAu151/ljg
By2m9or+S3rSy8gCat6zpoG4ZnLKJfonww3uOe/8fbbWG3zbRuWjQ+ufZn1hkFfx
15YCtzNorXReA4eSDpEX2rLBEOfTR2kB22YAV0aSxgMp7CD+HFdd7P/OwoMj7XWK
4HU/zMmU67yggaHHkZrnjL72kk7vzN4iqw3XhXgsTR/XgJd9Xhl8kXjZgCC2FpmZ
RyP6Ea4G5/tGl1F76Qh7gZEquQb7hIQXD2BRLyPSCzyXccCpcGYFc0/WPwehbKUQ
5g9KnEJVXhoPi/PFSW1GM/RccfzZsBo/vkVX8qt5RLIM20rgRD3hcfatA09Y6hsC
ryKD2Kpbf2PmzJCq/UlnDh9H7l7cDEvetSet4dYhJ2OVIy8OMvYdNAOBtBsnoOVY
zQbxxq818zzX+1CAyGGFd9j1jNtRTI7luxFRklFfkCG/kRqnyxvjvD+cViuaw4cO
mJnCGhNX5V8qkJ4vYrPblqYjetSZF3/EeZwR0KYte/qwaMROGId+2oMvQrQVMNmZ
L1GRm5eIlAPQOE5Qd09q/O9vljKt6FJQa8wP8DZ/Y1UukZbZ4ni/KieEKXp2Dsls
ouehGAwWNb98Kf/x2mTJEIIYcPBmmu3QC43cj2qZkSAZoLiyGiQZ5GU9+1ls4A5W
KF2VuYVku3cOjPjOcmFZ6JuLisZcBW2Y9IbmEnU60Vv2+kG48ZhwtJFvhBcQgqWu
Ns+sxwAJQ/7Zak7yIqc1Jx8bECDUdJTPI3cSh8eFc6vAe+jbRAvHhatxRRtArqxj
expk6/DLIjF6uGJ+5DHK4bb5NOaiI8gGiXYbAe6PUqK3R2BwvjJ/LJMgpmqUKMaj
dnnSLx1xsKCBPGmZjhgV6d1K+AzSHk2ZRZgTbUPt2DvoRXy4bFLNp/MPtcwz3Y9x
btmMdUHFMvupyPzU1hoQO+WWP3aystRSJ3YrRrHPD9AqUj4b3df1Qz/zycp1o6Sr
MJGjbTs8ziJP1cIhbrQpBU0tps5KsP1n7wp/mKaNdKTtYcZyScabMb7y74zFUYnb
yrKUk1eEdsXDvGTQnSQfr5p412EV4aVUwTEca3jVzUIE7nF7xTdUOKRHtG8nZJKd
7v0SNIHushHxPZh94wZKvNnNO7puKVtN3M7px/FBkZ3G1h2838vSd39tKIib1uUg
YrwLdZNW9uDjYVKYAYf+pkedkYNysByNKoHyNxD0lG6UHxX+h/JxSmWMkBQgRedS
6Rp0mxmJv4BvKIrEqHXM21giF7vBBnAB//ozHpg+xR7KRZbArMGnYCzO/mDyU8qr
TcQrsvmFqOE1C88aymBAJatHRuN/oh5RSAWO0umxLgnkImaXvgDvBzoA+G4/scsP
F5mKCKdtPWJ2J+z+TsXg8yF8YMDNdKaMsBaeeZVC2WlUsgpqB8VphaXfqRIBdpjX
fihbqDIcUrgeklS1D7FUXGAzH3mUWZ8CgrUCcDZ/HRtUSmdPREDeKp7ywbBYMpUw
9w2/tLGYyZVnGOB4nyVDssCd/qBdoI/Qa2FaQ0B+yzfQZpird/U5KBVOuXnMaRgi
2ML9TzoADlK+vuuqKjau2qdb8a22e7/rTSRYzzdbmNUQewFycuWPcEi7VLc8y+De
CUI03ybXS6kjrIShxw2qleRZDFto+sVJEQp/apBi480HNpULzE+BoKeGJPs4WvM1
WgtXdqTdqdJyvdC3hIr6QRwZQEzOP+que5iwBBM82fKPc7eKQjCXCNdFqoQ+WU4m
TJ5dBUUUg2CtT5dXKw3lpr0hTeDWhtkKqQbE3s1D4ZKYlC0yQ43wb1B2sjYGRghP
66ngRyqL+rk+vEv4ApTboSSLs6KCKqGqZEWhzJyDAP+c4Pe/fuhHOujX55kL1bUQ
jIQFFHtiaxLRO3WzjYVdfOCNfwDkNKCpHBFAtom/OmrrUqwC3MWy0Dv+IgNxETNo
Ihw3YSgu53v1l5HJTshCFj9af/lS2SSO5i1jyWQAOhNmuQxFfFWA73KlsrawtwXr
/8NF34KEbirXZnwvFKqIa9araciLhz2bmroys1Xl8ww529PiCk7axNXujn7nnLqO
ysZR3yr5BWkfpDQTykAzv7/EZmmJ1mdxkQ2DclkKQhTYrRBsERAP7Xk4CK2Bb7tA
2dR+K93fATpaVICEC9HoG8WWr3JH8FxIj1Un4IvxTPsLI6LT80zBq+AO1RYGMj4j
5B4w6uXVKm8Dpk79PqjTgz86/gCpxA++Vg2ReQcxX89788Kl5MT0kNuhQ0hBgABD
7mpHhcsG1zgOQ8f9n7Ci4fzpK4VJ6HacE2uo1KqYgVBxkyXgx3CJ/I/9i+jO7H3c
9w4cvzZ+VXb8D/auPaczPUsupUgZMaUT2WpHhNWppmGkRB4/d24E8mBmRkUPtuVx
IVlk/GOQMezUKsJ61l9o7xI0vnCGEFwCKaBmDOMIIggUf2bf34Pf0U6Le3pZ0nUW
hRyBVFNmLh/hLY+5wck4GGqNxNtGmNl1DlxIxig0M90BtwT9BSZyg/s96/aEeD33
xe+F86yr4hAMn5pZmysNfrjgq91/m84FhzCgW9X87O3umQfnwwV0IvVnYNVfRJfm
sIzLG3yvpsS2LJl/wRTUxl1xRwlPk/73rQ/G2B9oJ8HFFU/KGwheU+R/IA6RuCCP
p4jF0sfy1HGlD2EfYt0r4h5KS4PEv3Oo+eJg7MuqlREh2eylRG8bCw+DDVP3Q1SQ
b1MIlmHaOAfUFW3yet2MTouHVxNW+nsgRTxTkN6WkCm8QpXC+m6hMmt8fWzAIfOI
+6jsR1O5Klzk007B/4zaCcaOm/rTfDTiHNj7dmkemFfVvhgeHJqAVeZD7pMfV/x1
qRILGgLiZog89h/Q6cuylnPXhHz8MTehq2oWJfZdT7t4DgfvEnNZgdRVNpaHxTzr
ZS4+9J/foCUNlcQmc4ZLy/zgXQlLCsnhWjmCsqLt8imMvVi8peN5YycmCJfds5By
HJ+8B2mfsVPu1KCYmRVj/c7dTQeTZQC4LZi+Nl+WHSKBqVegBe0Oh0ot0xhBliej
9G9UvtUtRCL62/N4ISr15r6ERqhSblat76/h2vX5+PrftjlcPytLafLd8EaGOHxb
WqNEZgYkugU66eTYSPQ2/u+bi/n1XpknVN7imqBTVKO03kBPTMmG6dykpuy/8LyF
cVJFXvIgGj0HkB0Dm6EWTx4txliQ4M4yc+e7Eg1ctuUiI/RBsXzOv37rK8Vxy+F5
KOEbY2IFVlwS7VMNoyBrDZ52lBB1zbHif2fQxtcEsX6dJeB1MKHCve3JLyFSK8Qx
6+TuNeZTqcl1F1L7YpeRzGm2j2X6uoQEsaOLkatOWr5twnhaNZq6kmosgTeBeB/c
DAHVBsuKUypNuHsBP0OP8bl16CQb1p+dA8C9ZuX9CA3kd1374DdbS7tKnrVPScaU
YASuVWlVglOPJ/fX9FWRPs+g4W+yoqGvbpEZpie00in20ClKpVil7/p13dA+EkXN
myoCfDV5An82jE/lxilGnuIBr+Manz4j/0caOZyFeUvMwiwp3GcvvZ8k3CBFkK4E
Qh/Bx8ICQ60ZPqmOt/YCqNV4i0GbUOSEQiyb6LL+DcgoF7zdf5WqEurQ2AOG7j6d
atJkhRC+ZO7SC1yVAP9eT8wjHVH1jSFQmKYc363P+05WFxrTykilgAlg378qyEHF
Ir/umzy0JWDXqi6X/4+4Getb1Itt5m4aUbEIIhBBF6BDwazBwhjcDne65fXBJbI9
4eeYgiNzV8Z6raok6/yp1dfoI5+EuViEuXE0+m/ndTBtRD/vQnG3PshvNJ8joOcC
RGeE+38F48jsuV2bx8yvT+u7QWbQXTjrYFsrjJvL84pozg3y9v0wZ5eWQ3aZwRPs
n5zDKV/2oxrh2GlcYPfEkM0TGWZrreCEYVtNSvgZd19Hic8Kv/2S5CCdD3p2luMp
e+X/ifI4X+46JAYbWo1Yaz0uaqHlSd5ozi+iY45oEyO09ndIZo+R5unvAPZJqHfL
DjFOSCwG7dCxtCyx0xQT6X90HLDk/BIo4kRxHfI4I4pkpQz7XlZJNbQ/2vsaU31L
JtbOqHR0B4aHc+vi23jz4CXo2y+uIEutAsiklj45t0DLG6kGeIpYDkJVzx6PNN0Z
xeYSltElmQgN3oOveqfzGR3uunJUPUXwpTuVbzlq3D2twEzkpg7ZaZjLKOtzTGLM
R0tjACHWWsagOXJ/R7MKXGh6ir7XwUgFGLePlRBbGj0yhYcpWD/64oc/lfRbw1ev
u0HJ2L4Tl2fKlf41aduTNL2WpWxBd/VPpE4TSlYzw7zuDj1Y30WyCBQWVcTzXkkY
eLhBUr5tEqm2wXBzyKTUa9bd7CYTzdyuH3cwmcgn5dUGfMtXo1gB6YQNRhYSFEhJ
s22TUGRfeecGAbIV5FPljvp4fYlgjZJwo5vgg6Fw1v8JtIaM9+M/enSQ0Vhoky+d
vPzkQIJGCzcBjN+r9PNdNY1ItRtanCjMkrAW3f0I7+2azXE1vyRME0ibbdcmR5cz
PgSCZEEA7GTbFWngrlewrsaPqgHZUDqrs+wDdE+jiMCykr53CEhsXyQKtHod9Lid
OUucnrmydO0ynA0wpr3JReiNuYnLGsJK7thtqYi1QVfsSbS2fZVZ9wyxBtseiqV3
qp4VfbCM7+MtBozKQhdkfidbOHmHCgDtnhtQD/Tft2U=
`pragma protect end_protected
